
-- In this example, we're going to map voltage to distance, using a linear 
-- approximation, according to the Sharp GP2Y0A41SK0F datasheet page 4, or 
-- Lab 3 handout page 5. 
-- 
-- The relevant points we will select are:
-- 2.750 V is  4.00 cm (or 2750 mV and  40.0 mm)
-- 0.400 V is 33.00 cm (or  400 mV and 330.0 mm)
-- 
-- Mapping to the scales in our system
-- 2750 (mV) should map to  400 (10^-4 m)
--  400 (mV) should map to 3300 (10^-4 m)
-- and developing a linear equation, we find:
--
-- Distance = -2900/2350 * Voltage + 3793.617
-- Note this code implements linear function, you must map to the 
-- NON-linear relationship in the datasheet. This code is only provided 
-- for reference to help get you started.

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY BuzzFreq_Lookup IS
   PORT(
      clk            :  IN    STD_LOGIC;                                
      reset          :  IN    STD_LOGIC;                                
      index      	 :  IN    integer;                           
      Increment     :  OUT   integer
		);
END BuzzFreq_Lookup;

ARCHITECTURE behavior OF BuzzFreq_Lookup IS

type array_1d is array (0 to 4095) of Integer;

constant Increments : array_1d := (						
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(54975581),
(54976257),
(54976933),
(54977609),
(54978284),
(54978960),
(54979636),
(54980312),
(54980987),
(54981663),
(54982339),
(54983015),
(54983690),
(54984366),
(54985042),
(54985718),
(54986393),
(54987069),
(54987745),
(54988421),
(54989096),
(54989772),
(54990448),
(54991124),
(54991799),
(54992475),
(54993151),
(54993827),
(54994503),
(54995178),
(54995854),
(54996530),
(54997206),
(54997881),
(54998557),
(54999233),
(54999909),
(55000584),
(55001260),
(55001936),
(55002612),
(55003287),
(55003963),
(55004639),
(55005315),
(55005990),
(55006666),
(55007342),
(55008018),
(55008693),
(55009369),
(55010045),
(55010721),
(55011396),
(55012072),
(55012748),
(55013424),
(55014099),
(55014775),
(55015451),
(55016127),
(55016802),
(55017478),
(55018154),
(55018830),
(55019505),
(55020181),
(55020857),
(55021533),
(55022208),
(55022884),
(55023560),
(55024236),
(55024911),
(55025587),
(55026263),
(55026939),
(55027614),
(55028290),
(55028966),
(55029642),
(55030317),
(55030993),
(55031669),
(55032345),
(55033020),
(55033696),
(55034372),
(55035048),
(55035724),
(55036399),
(55037075),
(55037751),
(55038427),
(55039102),
(55039778),
(55040454),
(55041130),
(55041805),
(55042481),
(55043157),
(55043833),
(55044508),
(55045184),
(55045860),
(55046536),
(55047211),
(55047887),
(55048563),
(55049239),
(55049914),
(55050590),
(55051266),
(55051942),
(55052617),
(55053293),
(55053969),
(55054645),
(55055320),
(55055996),
(55056672),
(55057348),
(55058023),
(55058699),
(55059375),
(55060051),
(55060726),
(55061402),
(55062078),
(55062754),
(55063429),
(55064105),
(55064781),
(55065457),
(55066132),
(55066808),
(55067484),
(55068160),
(55068835),
(55069511),
(55070187),
(55070863),
(55071538),
(55072214),
(55072890),
(55073566),
(55074241),
(55074917),
(55075593),
(55076269),
(55076945),
(55077620),
(55078296),
(55078972),
(55079648),
(55080323),
(55080999),
(55081675),
(55082351),
(55083026),
(55083702),
(55084378),
(55085054),
(55085729),
(55086405),
(55087081),
(55087757),
(55088432),
(55089108),
(55089784),
(55090460),
(55091135),
(55091811),
(55092487),
(55093163),
(55093838),
(55094514),
(55095190),
(55095866),
(55096541),
(55097217),
(55097893),
(55098569),
(55099244),
(55099920),
(55100596),
(55101272),
(55101947),
(55102623),
(55103299),
(55103975),
(55104650),
(55105326),
(55106002),
(55106678),
(55107353),
(55108029),
(55108705),
(55109381),
(55110056),
(55110732),
(55111408),
(55112084),
(55112759),
(55113435),
(55114111),
(55114787),
(55115462),
(55116138),
(55116814),
(55117490),
(55118166),
(55118841),
(55119517),
(55120193),
(55120869),
(55121544),
(55122220),
(55122896),
(55123572),
(55124247),
(55124923),
(55125599),
(55126275),
(55126950),
(55127626),
(55128302),
(55128978),
(55129653),
(55130329),
(55131005),
(55131681),
(55132356),
(55133032),
(55133708),
(55134384),
(55135059),
(55135735),
(55136411),
(55137087),
(55137762),
(55138438),
(55139114),
(55139790),
(55140465),
(55141141),
(55141817),
(55142493),
(55143168),
(55143844),
(55144520),
(55145196),
(55145871),
(55146547),
(55147223),
(55147899),
(55148574),
(55149250),
(55149926),
(55150602),
(55151277),
(55151953),
(55152629),
(55153305),
(55153980),
(55154656),
(55155332),
(55156008),
(55156683),
(55157359),
(55158035),
(55158711),
(55159387),
(55160062),
(55160738),
(55161414),
(55162090),
(55162765),
(55163441),
(55164117),
(55164793),
(55165468),
(55166144),
(55166820),
(55167496),
(55168171),
(55168847),
(55169523),
(55170199),
(55170874),
(55171550),
(55172226),
(55172902),
(55173577),
(55174253),
(55174929),
(55175605),
(55176280),
(55176956),
(55177632),
(55178308),
(55178983),
(55179659),
(55180335),
(55181011),
(55181686),
(55182362),
(55183038),
(55183714),
(55184389),
(55185065),
(55185741),
(55186417),
(55187092),
(55187768),
(55188444),
(55189120),
(55189795),
(55190471),
(55191147),
(55191823),
(55192498),
(55193174),
(55193850),
(55194526),
(55195201),
(55195877),
(55196553),
(55197229),
(55197904),
(55198580),
(55199256),
(55199932),
(55200608),
(55201283),
(55201959),
(55202635),
(55203311),
(55203986),
(55204662),
(55205338),
(55206014),
(55206689),
(55207365),
(55208041),
(55208717),
(55209392),
(55210068),
(55210744),
(55211420),
(55212095),
(55212771),
(55213447),
(55214123),
(55214798),
(55215474),
(55216150),
(55216826),
(55217501),
(55218177),
(55218853),
(55219529),
(55220204),
(55220880),
(55221556),
(55222232),
(55222907),
(55223583),
(55224259),
(55224935),
(55225610),
(55226286),
(55226962),
(55227638),
(55228313),
(55228989),
(55229665),
(55230341),
(55231016),
(55231692),
(55232368),
(55233044),
(55233719),
(55234395),
(55235071),
(55235747),
(55236422),
(55237098),
(55237774),
(55238450),
(55239125),
(55239801),
(55240477),
(55241153),
(55241829),
(55242504),
(55243180),
(55243856),
(55244532),
(55245207),
(55245883),
(55246559),
(55247235),
(55247910),
(55248586),
(55249262),
(55249938),
(55250613),
(55251289),
(55251965),
(55252641),
(55253316),
(55253992),
(55254668),
(55255344),
(55256019),
(55256695),
(55257371),
(55258047),
(55258722),
(55259398),
(55260074),
(55260750),
(55261425),
(55262101),
(55262777),
(55263453),
(55264128),
(55264804),
(55265480),
(55266156),
(55266831),
(55267507),
(55268183),
(55268859),
(55269534),
(55270210),
(55270886),
(55271562),
(55272237),
(55272913),
(55273589),
(55274265),
(55274940),
(55275616),
(55276292),
(55276968),
(55277643),
(55278319),
(55278995),
(55279671),
(55280346),
(55281022),
(55281698),
(55282374),
(55283050),
(55283725),
(55284401),
(55285077),
(55285753),
(55286428),
(55287104),
(55287780),
(55288456),
(55289131),
(55289807),
(55290483),
(55291159),
(55291834),
(55292510),
(55293186),
(55293862),
(55294537),
(55295213),
(55295889),
(55296565),
(55297240),
(55297916),
(55298592),
(55299268),
(55299943),
(55300619),
(55301295),
(55301971),
(55302646),
(55303322),
(55303998),
(55304674),
(55305349),
(55306025),
(55306701),
(55307377),
(55308052),
(55308728),
(55309404),
(55310080),
(55310755),
(55311431),
(55312107),
(55312783),
(55313458),
(55314134),
(55314810),
(55315486),
(55316161),
(55316837),
(55317513),
(55318189),
(55318864),
(55319540),
(55320216),
(55320892),
(55321567),
(55322243),
(55322919),
(55323595),
(55324271),
(55324946),
(55325622),
(55326298),
(55326974),
(55327649),
(55328325),
(55329001),
(55329677),
(55330352),
(55331028),
(55331704),
(55332380),
(55333055),
(55333731),
(55334407),
(55335083),
(55335758),
(55336434),
(55337110),
(55337786),
(55338461),
(55339137),
(55339813),
(55340489),
(55341164),
(55341840),
(55342516),
(55343192),
(55343867),
(55344543),
(55345219),
(55345895),
(55346570),
(55347246),
(55347922),
(55348598),
(55349273),
(55349949),
(55350625),
(55351301),
(55351976),
(55352652),
(55353328),
(55354004),
(55354679),
(55355355),
(55356031),
(55356707),
(55357382),
(55358058),
(55358734),
(55359410),
(55360085),
(55360761),
(55361437),
(55362113),
(55362788),
(55363464),
(55364140),
(55364816),
(55365492),
(55366167),
(55366843),
(55367519),
(55368195),
(55368870),
(55369546),
(55370222),
(55370898),
(55371573),
(55372249),
(55372925),
(55373601),
(55374276),
(55374952),
(55375628),
(55376304),
(55376979),
(55377655),
(55378331),
(55379007),
(55379682),
(55380358),
(55381034),
(55381710),
(55382385),
(55383061),
(55383737),
(55384413),
(55385088),
(55385764),
(55386440),
(55387116),
(55387791),
(55388467),
(55389143),
(55389819),
(55390494),
(55391170),
(55391846),
(55392522),
(55393197),
(55393873),
(55394549),
(55395225),
(55395900),
(55396576),
(55397252),
(55397928),
(55398603),
(55399279),
(55399955),
(55400631),
(55401306),
(55401982),
(55402658),
(55403334),
(55404009),
(55404685),
(55405361),
(55406037),
(55406713),
(55407388),
(55408064),
(55408740),
(55409416),
(55410091),
(55410767),
(55411443),
(55412119),
(55412794),
(55413470),
(55414146),
(55414822),
(55415497),
(55416173),
(55416849),
(55417525),
(55418200),
(55418876),
(55419552),
(55420228),
(55420903),
(55421579),
(55422255),
(55422931),
(55423606),
(55424282),
(55424958),
(55425634),
(55426309),
(55426985),
(55427661),
(55428337),
(55429012),
(55429688),
(55430364),
(55431040),
(55431715),
(55432391),
(55433067),
(55433743),
(55434418),
(55435094),
(55435770),
(55436446),
(55437121),
(55437797),
(55438473),
(55439149),
(55439824),
(55440500),
(55441176),
(55441852),
(55442527),
(55443203),
(55443879),
(55444555),
(55445230),
(55445906),
(55446582),
(55447258),
(55447934),
(55448609),
(55449285),
(55449961),
(55450637),
(55451312),
(55451988),
(55452664),
(55453340),
(55454015),
(55454691),
(55455367),
(55456043),
(55456718),
(55457394),
(55458070),
(55458746),
(55459421),
(55460097),
(55460773),
(55461449),
(55462124),
(55462800),
(55463476),
(55464152),
(55464827),
(55465503),
(55466179),
(55466855),
(55467530),
(55468206),
(55468882),
(55469558),
(55470233),
(55470909),
(55471585),
(55472261),
(55472936),
(55473612),
(55474288),
(55474964),
(55475639),
(55476315),
(55476991),
(55477667),
(55478342),
(55479018),
(55479694),
(55480370),
(55481045),
(55481721),
(55482397),
(55483073),
(55483748),
(55484424),
(55485100),
(55485776),
(55486451),
(55487127),
(55487803),
(55488479),
(55489154),
(55489830),
(55490506),
(55491182),
(55491858),
(55492533),
(55493209),
(55493885),
(55494561),
(55495236),
(55495912),
(55496588),
(55497264),
(55497939),
(55498615),
(55499291),
(55499967),
(55500642),
(55501318),
(55501994),
(55502670),
(55503345),
(55504021),
(55504697),
(55505373),
(55506048),
(55506724),
(55507400),
(55508076),
(55508751),
(55509427),
(55510103),
(55510779),
(55511454),
(55512130),
(55512806),
(55513482),
(55514157),
(55514833),
(55515509),
(55516185),
(55516860),
(55517536),
(55518212),
(55518888),
(55519563),
(55520239),
(55520915),
(55521591),
(55522266),
(55522942),
(55523618),
(55524294),
(55524969),
(55525645),
(55526321),
(55526997),
(55527672),
(55528348),
(55529024),
(55529700),
(55530375),
(55531051),
(55531727),
(55532403),
(55533079),
(55533754),
(55534430),
(55535106),
(55535782),
(55536457),
(55537133),
(55537809),
(55538485),
(55539160),
(55539836),
(55540512),
(55541188),
(55541863),
(55542539),
(55543215),
(55543891),
(55544566),
(55545242),
(55545918),
(55546594),
(55547269),
(55547945),
(55548621),
(55549297),
(55549972),
(55550648),
(55551324),
(55552000),
(55552675),
(55553351),
(55554027),
(55554703),
(55555378),
(55556054),
(55556730),
(55557406),
(55558081),
(55558757),
(55559433),
(55560109),
(55560784),
(55561460),
(55562136),
(55562812),
(55563487),
(55564163),
(55564839),
(55565515),
(55566190),
(55566866),
(55567542),
(55568218),
(55568893),
(55569569),
(55570245),
(55570921),
(55571596),
(55572272),
(55572948),
(55573624),
(55574300),
(55574975),
(55575651),
(55576327),
(55577003),
(55577678),
(55578354),
(55579030),
(55579706),
(55580381),
(55581057),
(55581733),
(55582409),
(55583084),
(55583760),
(55584436),
(55585112),
(55585787),
(55586463),
(55587139),
(55587815),
(55588490),
(55589166),
(55589842),
(55590518),
(55591193),
(55591869),
(55592545),
(55593221),
(55593896),
(55594572),
(55595248),
(55595924),
(55596599),
(55597275),
(55597951),
(55598627),
(55599302),
(55599978),
(55600654),
(55601330),
(55602005),
(55602681),
(55603357),
(55604033),
(55604708),
(55605384),
(55606060),
(55606736),
(55607411),
(55608087),
(55608763),
(55609439),
(55610114),
(55610790),
(55611466),
(55612142),
(55612817),
(55613493),
(55614169),
(55614845),
(55615521),
(55616196),
(55616872),
(55617548),
(55618224),
(55618899),
(55619575),
(55620251),
(55620927),
(55621602),
(55622278),
(55622954),
(55623630),
(55624305),
(55624981),
(55625657),
(55626333),
(55627008),
(55627684),
(55628360),
(55629036),
(55629711),
(55630387),
(55631063),
(55631739),
(55632414),
(55633090),
(55633766),
(55634442),
(55635117),
(55635793),
(55636469),
(55637145),
(55637820),
(55638496),
(55639172),
(55639848),
(55640523),
(55641199),
(55641875),
(55642551),
(55643226),
(55643902),
(55644578),
(55645254),
(55645929),
(55646605),
(55647281),
(55647957),
(55648632),
(55649308),
(55649984),
(55650660),
(55651335),
(55652011),
(55652687),
(55653363),
(55654038),
(55654714),
(55655390),
(55656066),
(55656742),
(55657417),
(55658093),
(55658769),
(55659445),
(55660120),
(55660796),
(55661472),
(55662148),
(55662823),
(55663499),
(55664175),
(55664851),
(55665526),
(55666202),
(55666878),
(55667554),
(55668229),
(55668905),
(55669581),
(55670257),
(55670932),
(55671608),
(55672284),
(55672960),
(55673635),
(55674311),
(55674987),
(55675663),
(55676338),
(55677014),
(55677690),
(55678366),
(55679041),
(55679717),
(55680393),
(55681069),
(55681744),
(55682420),
(55683096),
(55683772),
(55684447),
(55685123),
(55685799),
(55686475),
(55687150),
(55687826),
(55688502),
(55689178),
(55689853),
(55690529),
(55691205),
(55691881),
(55692556),
(55693232),
(55693908),
(55694584),
(55695259),
(55695935),
(55696611),
(55697287),
(55697963),
(55698638),
(55699314),
(55699990),
(55700666),
(55701341),
(55702017),
(55702693),
(55703369),
(55704044),
(55704720),
(55705396),
(55706072),
(55706747),
(55707423),
(55708099),
(55708775),
(55709450),
(55710126),
(55710802),
(55711478),
(55712153),
(55712829),
(55713505),
(55714181),
(55714856),
(55715532),
(55716208),
(55716884),
(55717559),
(55718235),
(55718911),
(55719587),
(55720262),
(55720938),
(55721614),
(55722290),
(55722965),
(55723641),
(55724317),
(55724993),
(55725668),
(55726344),
(55727020),
(55727696),
(55728371),
(55729047),
(55729723),
(55730399),
(55731074),
(55731750),
(55732426),
(55733102),
(55733777),
(55734453),
(55735129),
(55735805),
(55736480),
(55737156),
(55737832),
(55738508),
(55739184),
(55739859),
(55740535),
(55741211),
(55741887),
(55742562),
(55743238),
(55743914),
(55744590),
(55745265),
(55745941),
(55746617),
(55747293),
(55747968),
(55748644),
(55749320),
(55749996),
(55750671),
(55751347),
(55752023),
(55752699),
(55753374),
(55754050),
(55754726),
(55755402),
(55756077),
(55756753),
(55757429),
(55758105),
(55758780),
(55759456),
(55760132),
(55760808),
(55761483),
(55762159),
(55762835),
(55763511),
(55764186),
(55764862),
(55765538),
(55766214),
(55766889),
(55767565),
(55768241),
(55768917),
(55769592),
(55770268),
(55770944),
(55771620),
(55772295),
(55772971),
(55773647),
(55774323),
(55774998),
(55775674),
(55776350),
(55777026),
(55777701),
(55778377),
(55779053),
(55779729),
(55780405),
(55781080),
(55781756),
(55782432),
(55783108),
(55783783),
(55784459),
(55785135),
(55785811),
(55786486),
(55787162),
(55787838),
(55788514),
(55789189),
(55789865),
(55790541),
(55791217),
(55791892),
(55792568),
(55793244),
(55793920),
(55794595),
(55795271),
(55795947),
(55796623),
(55797298),
(55797974),
(55798650),
(55799326),
(55800001),
(55800677),
(55801353),
(55802029),
(55802704),
(55803380),
(55804056),
(55804732),
(55805407),
(55806083),
(55806759),
(55807435),
(55808110),
(55808786),
(55809462),
(55810138),
(55810813),
(55811489),
(55812165),
(55812841),
(55813516),
(55814192),
(55814868),
(55815544),
(55816219),
(55816895),
(55817571),
(55818247),
(55818922),
(55819598),
(55820274),
(55820950),
(55821626),
(55822301),
(55822977),
(55823653),
(55824329),
(55825004),
(55825680),
(55826356),
(55827032),
(55827707),
(55828383),
(55829059),
(55829735),
(55830410),
(55831086),
(55831762),
(55832438),
(55833113),
(55833789),
(55834465),
(55835141),
(55835816),
(55836492),
(55837168),
(55837844),
(55838519),
(55839195),
(55839871),
(55840547),
(55841222),
(55841898),
(55842574),
(55843250),
(55843925),
(55844601),
(55845277),
(55845953),
(55846628),
(55847304),
(55847980),
(55848656),
(55849331),
(55850007),
(55850683),
(55851359),
(55852034),
(55852710),
(55853386),
(55854062),
(55854737),
(55855413),
(55856089),
(55856765),
(55857440),
(55858116),
(55858792),
(55859468),
(55860143),
(55860819),
(55861495),
(55862171),
(55862847),
(55863522),
(55864198),
(55864874),
(55865550),
(55866225),
(55866901),
(55867577),
(55868253),
(55868928),
(55869604),
(55870280),
(55870956),
(55871631),
(55872307),
(55872983),
(55873659),
(55874334),
(55875010),
(55875686),
(55876362),
(55877037),
(55877713),
(55878389),
(55879065),
(55879740),
(55880416),
(55881092),
(55881768),
(55882443),
(55883119),
(55883795),
(55884471),
(55885146),
(55885822),
(55886498),
(55887174),
(55887849),
(55888525),
(55889201),
(55889877),
(55890552),
(55891228),
(55891904),
(55892580),
(55893255),
(55893931),
(55894607),
(55895283),
(55895958),
(55896634),
(55897310),
(55897986),
(55898661),
(55899337),
(55900013),
(55900689),
(55901364),
(55902040),
(55902716),
(55903392),
(55904068),
(55904743),
(55905419),
(55906095),
(55906771),
(55907446),
(55908122),
(55908798),
(55909474),
(55910149),
(55910825),
(55911501),
(55912177),
(55912852),
(55913528),
(55914204),
(55914880),
(55915555),
(55916231),
(55916907),
(55917583),
(55918258),
(55918934),
(55919610),
(55920286),
(55920961),
(55921637),
(55922313),
(55922989),
(55923664),
(55924340),
(55925016),
(55925692),
(55926367),
(55927043),
(55927719),
(55928395),
(55929070),
(55929746),
(55930422),
(55931098),
(55931773),
(55932449),
(55933125),
(55933801),
(55934476),
(55935152),
(55935828),
(55936504),
(55937179),
(55937855),
(55938531),
(55939207),
(55939882),
(55940558),
(55941234),
(55941910),
(55942585),
(55943261),
(55943937),
(55944613),
(55945289),
(55945964),
(55946640),
(55947316),
(55947992),
(55948667),
(55949343),
(55950019),
(55950695),
(55951370),
(55952046),
(55952722),
(55953398),
(55954073),
(55954749),
(55955425),
(55956101),
(55956776),
(55957452),
(55958128),
(55958804),
(55959479),
(55960155),
(55960831),
(55961507),
(55962182),
(55962858),
(55963534),
(55964210),
(55964885),
(55965561),
(55966237),
(55966913),
(55967588),
(55968264),
(55968940),
(55969616),
(55970291),
(55970967),
(55971643),
(55972319),
(55972994),
(55973670),
(55974346),
(55975022),
(55975697),
(55976373),
(55977049),
(55977725),
(55978400),
(55979076),
(55979752),
(55980428),
(55981103),
(55981779),
(55982455),
(55983131),
(55983806),
(55984482),
(55985158),
(55985834),
(55986510),
(55987185),
(55987861),
(55988537),
(55989213),
(55989888),
(55990564),
(55991240),
(55991916),
(55992591),
(55993267),
(55993943),
(55994619),
(55995294),
(55995970),
(55996646),
(55997322),
(55997997),
(55998673),
(55999349),
(56000025),
(56000700),
(56001376),
(56002052),
(56002728),
(56003403),
(56004079),
(56004755),
(56005431),
(56006106),
(56006782),
(56007458),
(56008134),
(56008809),
(56009485),
(56010161),
(56010837),
(56011512),
(56012188),
(56012864),
(56013540),
(56014215),
(56014891),
(56015567),
(56016243),
(56016918),
(56017594),
(56018270),
(56018946),
(56019621),
(56020297),
(56020973),
(56021649),
(56022324),
(56023000),
(56023676),
(56024352),
(56025027),
(56025703),
(56026379),
(56027055),
(56027731),
(56028406),
(56029082),
(56029758),
(56030434),
(56031109),
(56031785),
(56032461),
(56033137),
(56033812),
(56034488),
(56035164),
(56035840),
(56036515),
(56037191),
(56037867),
(56038543),
(56039218),
(56039894),
(56040570),
(56041246),
(56041921),
(56042597),
(56043273),
(56043949),
(56044624),
(56045300),
(56045976),
(56046652),
(56047327),
(56048003),
(56048679),
(56049355),
(56050030),
(56050706),
(56051382),
(56052058),
(56052733),
(56053409),
(56054085),
(56054761),
(56055436),
(56056112),
(56056788),
(56057464),
(56058139),
(56058815),
(56059491),
(56060167),
(56060842),
(56061518),
(56062194),
(56062870),
(56063545),
(56064221),
(56064897),
(56065573),
(56066248),
(56066924),
(56067600),
(56068276),
(56068952),
(56069627),
(56070303),
(56070979),
(56071655),
(56072330),
(56073006),
(56073682),
(56074358),
(56075033),
(56075709),
(56076385),
(56077061),
(56077736),
(56078412),
(56079088),
(56079764),
(56080439),
(56081115),
(56081791),
(56082467),
(56083142),
(56083818),
(56084494),
(56085170),
(56085845),
(56086521),
(56087197),
(56087873),
(56088548),
(56089224),
(56089900),
(56090576),
(56091251),
(56091927),
(56092603),
(56093279),
(56093954),
(56094630),
(56095306),
(56095982),
(56096657),
(56097333),
(56098009),
(56098685),
(56099360),
(56100036),
(56100712),
(56101388),
(56102063),
(56102739),
(56103415),
(56104091),
(56104766),
(56105442),
(56106118),
(56106794),
(56107469),
(56108145),
(56108821),
(56109497),
(56110173),
(56110848),
(56111524),
(56112200),
(56112876),
(56113551),
(56114227),
(56114903),
(56115579),
(56116254),
(56116930),
(56117606),
(56118282),
(56118957),
(56119633),
(56120309),
(56120985),
(56121660),
(56122336),
(56123012),
(56123688),
(56124363),
(56125039),
(56125715),
(56126391),
(56127066),
(56127742),
(56128418),
(56129094),
(56129769),
(56130445),
(56131121),
(56131797),
(56132472),
(56133148),
(56133824),
(56134500),
(56135175),
(56135851),
(56136527),
(56137203),
(56137878),
(56138554),
(56139230),
(56139906),
(56140581),
(56141257),
(56141933),
(56142609),
(56143284),
(56143960),
(56144636),
(56145312),
(56145987),
(56146663),
(56147339),
(56148015),
(56148690),
(56149366),
(56150042),
(56150718),
(56151394),
(56152069),
(56152745),
(56153421),
(56154097),
(56154772),
(56155448),
(56156124),
(56156800),
(56157475),
(56158151),
(56158827),
(56159503),
(56160178),
(56160854),
(56161530),
(56162206),
(56162881),
(56163557),
(56164233),
(56164909),
(56165584),
(56166260),
(56166936),
(56167612),
(56168287),
(56168963),
(56169639),
(56170315),
(56170990),
(56171666),
(56172342),
(56173018),
(56173693),
(56174369),
(56175045),
(56175721),
(56176396),
(56177072),
(56177748),
(56178424),
(56179099),
(56179775),
(56180451),
(56181127),
(56181802),
(56182478),
(56183154),
(56183830),
(56184505),
(56185181),
(56185857),
(56186533),
(56187208),
(56187884),
(56188560),
(56189236),
(56189911),
(56190587),
(56191263),
(56191939),
(56192615),
(56193290),
(56193966),
(56194642),
(56195318),
(56195993),
(56196669),
(56197345),
(56198021),
(56198696),
(56199372),
(56200048),
(56200724),
(56201399),
(56202075),
(56202751),
(56203427),
(56204102),
(56204778),
(56205454),
(56206130),
(56206805),
(56207481),
(56208157),
(56208833),
(56209508),
(56210184),
(56210860),
(56211536),
(56212211),
(56212887),
(56213563),
(56214239),
(56214914),
(56215590),
(56216266),
(56216942),
(56217617),
(56218293),
(56218969),
(56219645),
(56220320),
(56220996),
(56221672),
(56222348),
(56223023),
(56223699),
(56224375),
(56225051),
(56225726),
(56226402),
(56227078),
(56227754),
(56228429),
(56229105),
(56229781),
(56230457),
(56231132),
(56231808),
(56232484),
(56233160),
(56233836),
(56234511),
(56235187),
(56235863),
(56236539),
(56237214),
(56237890),
(56238566),
(56239242),
(56239917),
(56240593),
(56241269),
(56241945),
(56242620),
(56243296),
(56243972),
(56244648),
(56245323),
(56245999),
(56246675),
(56247351),
(56248026),
(56248702),
(56249378),
(56250054),
(56250729),
(56251405),
(56252081),
(56252757),
(56253432),
(56254108),
(56254784),
(56255460),
(56256135),
(56256811),
(56257487),
(56258163),
(56258838),
(56259514),
(56260190),
(56260866),
(56261541),
(56262217),
(56262893),
(56263569),
(56264244),
(56264920),
(56265596),
(56266272),
(56266947),
(56267623),
(56268299),
(56268975),
(56269650),
(56270326),
(56271002),
(56271678),
(56272353),
(56273029),
(56273705),
(56274381),
(56275057),
(56275732),
(56276408),
(56277084),
(56277760),
(56278435),
(56279111),
(56279787),
(56280463),
(56281138),
(56281814),
(56282490),
(56283166),
(56283841),
(56284517),
(56285193),
(56285869),
(56286544),
(56287220),
(56287896),
(56288572),
(56289247),
(56289923),
(56290599),
(56291275),
(56291950),
(56292626),
(56293302),
(56293978),
(56294653),
(56295329),
(56296005),
(56296681),
(56297356),
(56298032),
(56298708),
(56299384),
(56300059),
(56300735),
(56301411),
(56302087),
(56302762),
(56303438),
(56304114),
(56304790),
(56305465),
(56306141),
(56306817),
(56307493),
(56308168),
(56308844),
(56309520),
(56310196),
(56310871),
(56311547),
(56312223),
(56312899),
(56313574),
(56314250),
(56314926),
(56315602),
(56316278),
(56316953),
(56317629),
(56318305),
(56318981),
(56319656),
(56320332),
(56321008),
(56321684),
(56322359),
(56323035),
(56323711),
(56324387),
(56325062),
(56325738),
(56326414),
(56327090),
(56327765),
(56328441),
(56329117),
(56329793),
(56330468),
(56331144),
(56331820),
(56332496),
(56333171),
(56333847),
(56334523),
(56335199),
(56335874),
(56336550),
(56337226),
(56337902),
(56338577),
(56339253),
(56339929),
(56340605),
(56341280),
(56341956),
(56342632),
(56343308),
(56343983),
(56344659),
(56345335),
(56346011),
(56346686),
(56347362),
(56348038),
(56348714),
(56349389),
(56350065),
(56350741),
(56351417),
(56352092),
(56352768),
(56353444),
(56354120),
(56354795),
(56355471),
(56356147),
(56356823),
(56357499),
(56358174),
(56358850),
(56359526),
(56360202),
(56360877),
(56361553),
(56362229),
(56362905),
(56363580),
(56364256),
(56364932),
(56365608),
(56366283),
(56366959),
(56367635),
(56368311),
(56368986),
(56369662),
(56370338),
(56371014),
(56371689),
(56372365),
(56373041),
(56373717),
(56374392),
(56375068),
(56375744),
(56376420),
(56377095),
(56377771),
(56378447),
(56379123),
(56379798),
(56380474),
(56381150),
(56381826),
(56382501),
(56383177),
(56383853),
(56384529),
(56385204),
(56385880),
(56386556),
(56387232),
(56387907),
(56388583),
(56389259),
(56389935),
(56390610),
(56391286),
(56391962),
(56392638),
(56393313),
(56393989),
(56394665),
(56395341),
(56396016),
(56396692),
(56397368),
(56398044),
(56398720),
(56399395),
(56400071),
(56400747),
(56401423),
(56402098),
(56402774),
(56403450),
(56404126),
(56404801),
(56405477),
(56406153),
(56406829),
(56407504),
(56408180),
(56408856),
(56409532),
(56410207),
(56410883),
(56411559),
(56412235),
(56412910),
(56413586),
(56414262),
(56414938),
(56415613),
(56416289),
(56416965),
(56417641),
(56418316),
(56418992),
(56419668),
(56420344),
(56421019),
(56421695),
(56422371),
(56423047),
(56423722),
(56424398),
(56425074),
(56425750),
(56426425),
(56427101),
(56427777),
(56428453),
(56429128),
(56429804),
(56430480),
(56431156),
(56431831),
(56432507),
(56433183),
(56433859),
(56434534),
(56435210),
(56435886),
(56436562),
(56437237),
(56437913),
(56438589),
(56439265),
(56439941),
(56440616),
(56441292),
(56441968),
(56442644),
(56443319),
(56443995),
(56444671),
(56445347),
(56446022),
(56446698),
(56447374),
(56448050),
(56448725),
(56449401),
(56450077),
(56450753),
(56451428),
(56452104),
(56452780),
(56453456),
(56454131),
(56454807),
(56455483),
(56456159),
(56456834),
(56457510),
(56458186),
(56458862),
(56459537),
(56460213),
(56460889),
(56461565),
(56462240),
(56462916),
(56463592),
(56464268),
(56464943),
(56465619),
(56466295),
(56466971),
(56467646),
(56468322),
(56468998),
(56469674),
(56470349),
(56471025),
(56471701),
(56472377),
(56473052),
(56473728),
(56474404),
(56475080),
(56475755),
(56476431),
(56477107),
(56477783),
(56478458),
(56479134),
(56479810),
(56480486),
(56481162),
(56481837),
(56482513),
(56483189),
(56483865),
(56484540),
(56485216),
(56485892),
(56486568),
(56487243),
(56487919),
(56488595),
(56489271),
(56489946),
(56490622),
(56491298),
(56491974),
(56492649),
(56493325),
(56494001),
(56494677),
(56495352),
(56496028),
(56496704),
(56497380),
(56498055),
(56498731),
(56499407),
(56500083),
(56500758),
(56501434),
(56502110),
(56502786),
(56503461),
(56504137),
(56504813),
(56505489),
(56506164),
(56506840),
(56507516),
(56508192),
(56508867),
(56509543),
(56510219),
(56510895),
(56511570),
(56512246),
(56512922),
(56513598),
(56514273),
(56514949),
(56515625),
(56516301),
(56516976),
(56517652),
(56518328),
(56519004),
(56519679),
(56520355),
(56521031),
(56521707),
(56522383),
(56523058),
(56523734),
(56524410),
(56525086),
(56525761),
(56526437),
(56527113),
(56527789),
(56528464),
(56529140),
(56529816),
(56530492),
(56531167),
(56531843),
(56532519),
(56533195),
(56533870),
(56534546),
(56535222),
(56535898),
(56536573),
(56537249),
(56537925),
(56538601),
(56539276),
(56539952),
(56540628),
(56541304),
(56541979),
(56542655),
(56543331),
(56544007),
(56544682),
(56545358),
(56546034),
(56546710),
(56547385),
(56548061),
(56548737),
(56549413),
(56550088),
(56550764),
(56551440),
(56552116),
(56552791),
(56553467),
(56554143),
(56554819),
(56555494),
(56556170),
(56556846),
(56557522),
(56558197),
(56558873),
(56559549),
(56560225),
(56560900),
(56561576),
(56562252),
(56562928),
(56563604),
(56564279),
(56564955),
(56565631),
(56566307),
(56566982),
(56567658),
(56568334),
(56569010),
(56569685),
(56570361),
(56571037),
(56571713),
(56572388),
(56573064),
(56573740),
(56574416),
(56575091),
(56575767),
(56576443),
(56577119),
(56577794),
(56578470),
(56579146),
(56579822),
(56580497),
(56581173),
(56581849),
(56582525),
(56583200),
(56583876),
(56584552),
(56585228),
(56585903),
(56586579),
(56587255),
(56587931),
(56588606),
(56589282),
(56589958),
(56590634),
(56591309),
(56591985),
(56592661),
(56593337),
(56594012),
(56594688),
(56595364),
(56596040),
(56596715),
(56597391),
(56598067),
(56598743),
(56599418),
(56600094),
(56600770),
(56601446),
(56602121),
(56602797),
(56603473),
(56604149),
(56604825),
(56605500),
(56606176),
(56606852),
(56607528),
(56608203),
(56608879),
(56609555),
(56610231),
(56610906),
(56611582),
(56612258),
(56612934),
(56613609),
(56614285),
(56614961),
(56615637),
(56616312),
(56616988),
(56617664),
(56618340),
(56619015),
(56619691),
(56620367),
(56621043),
(56621718),
(56622394),
(56623070),
(56623746),
(56624421),
(56625097),
(56625773),
(56626449),
(56627124),
(56627800),
(56628476),
(56629152),
(56629827),
(56630503),
(56631179),
(56631855),
(56632530),
(56633206),
(56633882),
(56634558),
(56635233),
(56635909),
(56636585),
(56637261),
(56637936),
(56638612),
(56639288),
(56639964),
(56640639),
(56641315),
(56641991),
(56642667),
(56643342),
(56644018),
(56644694),
(56645370),
(56646046),
(56646721),
(56647397),
(56648073),
(56648749),
(56649424),
(56650100),
(56650776),
(56651452),
(56652127),
(56652803),
(56653479),
(56654155),
(56654830),
(56655506),
(56656182),
(56656858),
(56657533),
(56658209),
(56658885),
(56659561),
(56660236),
(56660912),
(56661588),
(56662264),
(56662939),
(56663615),
(56664291),
(56664967),
(56665642),
(56666318),
(56666994),
(56667670),
(56668345),
(56669021),
(56669697),
(56670373),
(56671048),
(56671724),
(56672400),
(56673076),
(56673751),
(56674427),
(56675103),
(56675779),
(56676454),
(56677130),
(56677806),
(56678482),
(56679157),
(56679833),
(56680509),
(56681185),
(56681860),
(56682536),
(56683212),
(56683888),
(56684563),
(56685239),
(56685915),
(56686591),
(56687267),
(56687942),
(56688618),
(56689294),
(56689970),
(56690645),
(56691321),
(56691997),
(56692673),
(56693348),
(56694024),
(56694700),
(56695376),
(56696051),
(56696727),
(56697403),
(56698079),
(56698754),
(56699430),
(56700106),
(56700782),
(56701457),
(56702133),
(56702809),
(56703485),
(56704160),
(56704836),
(56705512),
(56706188),
(56706863),
(56707539),
(56708215),
(56708891),
(56709566),
(56710242),
(56710918),
(56711594),
(56712269),
(56712945),
(56713621),
(56714297),
(56714972),
(56715648),
(56716324),
(56717000),
(56717675),
(56718351),
(56719027),
(56719703),
(56720378),
(56721054),
(56721730),
(56722406),
(56723081),
(56723757),
(56724433),
(56725109),
(56725784),
(56726460),
(56727136),
(56727812),
(56728488),
(56729163),
(56729839),
(56730515),
(56731191),
(56731866),
(56732542),
(56733218),
(56733894),
(56734569),
(56735245),
(56735921),
(56736597),
(56737272),
(56737948),
(56738624),
(56739300),
(56739975),
(56740651),
(56741327),
(56742003),
(56742678),
(56743354),
(56744030),
(56744706),
(56745381),
(56746057),
(56746733),
(56747409),
(56748084),
(56748760),
(56749436),
(56750112),
(56750787),
(56751463),
(56752139),
(56752815),
(56753490),
(56754166),
(56754842),
(56755518),
(56756193),
(56756869),
(56757545),
(56758221),
(56758896),
(56759572),
(56760248),
(56760924),
(56761599),
(56762275),
(56762951),
(56763627),
(56764302),
(56764978),
(56765654),
(56766330),
(56767005),
(56767681),
(56768357),
(56769033),
(56769709),
(56770384),
(56771060),
(56771736),
(56772412),
(56773087),
(56773763),
(56774439),
(56775115),
(56775790),
(56776466),
(56777142),
(56777818),
(56778493),
(56779169),
(56779845),
(56780521),
(56781196),
(56781872),
(56782548),
(56783224),
(56783899),
(56784575),
(56785251),
(56785927),
(56786602),
(56787278),
(56787954),
(56788630),
(56789305),
(56789981),
(56790657),
(56791333),
(56792008),
(56792684),
(56793360),
(56794036),
(56794711),
(56795387),
(56796063),
(56796739),
(56797414),
(56798090),
(56798766),
(56799442),
(56800117),
(56800793),
(56801469),
(56802145),
(56802820),
(56803496),
(56804172),
(56804848),
(56805523),
(56806199),
(56806875),
(56807551),
(56808226),
(56808902),
(56809578),
(56810254),
(56810930),
(56811605),
(56812281),
(56812957),
(56813633),
(56814308),
(56814984),
(56815660),
(56816336),
(56817011),
(56817687),
(56818363),
(56819039),
(56819714),
(56820390),
(56821066),
(56821742),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575)
);


begin
    -- This is the only statement required. It looks up the converted value of 
	-- the voltage input (in mV) in the v2d_LUT look-up table, and outputs the 
	-- distance (in 10^-4 m) in std_logic_vector format.
	yeet : process(index)
	begin
		if(index < 0) then
			Increment <= 55834575;
		elsif (index > 4095) then
			Increment <= 55834575;
		else
			Increment <= Increments(index);
		end if;
	end process;
--   distance <= std_logic_vector(to_unsigned(v2d_LUTshort(to_integer(unsigned(voltage))),distance'length));
--   distance <= std_logic_vector(to_unsigned(v2d_LUT(to_integer(unsigned(voltage))),distance'length));

end behavior;
