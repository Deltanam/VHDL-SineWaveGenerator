
-- In this example, we're going to map voltage to distance, using a linear 
-- approximation, according to the Sharp GP2Y0A41SK0F datasheet page 4, or 
-- Lab 3 handout page 5. 
-- 
-- The relevant points we will select are:
-- 2.750 V is  4.00 cm (or 2750 mV and  40.0 mm)
-- 0.400 V is 33.00 cm (or  400 mV and 330.0 mm)
-- 
-- Mapping to the scales in our system
-- 2750 (mV) should map to  400 (10^-4 m)
--  400 (mV) should map to 3300 (10^-4 m)
-- and developing a linear equation, we find:
--
-- Distance = -2900/2350 * Voltage + 3793.617
-- Note this code implements linear function, you must map to the 
-- NON-linear relationship in the datasheet. This code is only provided 
-- for reference to help get you started.

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY Sine_Lookup IS
   PORT(
      clk            :  IN    STD_LOGIC;                                
      reset          :  IN    STD_LOGIC;                                
      index      	 	:  IN    integer;                           
      duty_cycle     :  OUT   STD_LOGIC_VECTOR(9 downto 0)
		);
END Sine_Lookup;

ARCHITECTURE behavior OF Sine_Lookup IS

type array_1d is array (0 to 1023) of STD_LOGIC_VECTOR(9 downto 0);

constant Sinevalues : array_1d := (												
(	"0111111111"	)	,
(	"1000000010"	)	,
(	"1000000101"	)	,
(	"1000001000"	)	,
(	"1000001011"	)	,
(	"1000001110"	)	,
(	"1000010001"	)	,
(	"1000010100"	)	,
(	"1000011000"	)	,
(	"1000011011"	)	,
(	"1000011110"	)	,
(	"1000100001"	)	,
(	"1000100100"	)	,
(	"1000100111"	)	,
(	"1000101010"	)	,
(	"1000101101"	)	,
(	"1000110001"	)	,
(	"1000110100"	)	,
(	"1000110111"	)	,
(	"1000111010"	)	,
(	"1000111101"	)	,
(	"1001000000"	)	,
(	"1001000011"	)	,
(	"1001000110"	)	,
(	"1001001001"	)	,
(	"1001001101"	)	,
(	"1001010000"	)	,
(	"1001010011"	)	,
(	"1001010110"	)	,
(	"1001011001"	)	,
(	"1001011100"	)	,
(	"1001011111"	)	,
(	"1001100010"	)	,
(	"1001100101"	)	,
(	"1001101000"	)	,
(	"1001101011"	)	,
(	"1001101110"	)	,
(	"1001110010"	)	,
(	"1001110101"	)	,
(	"1001111000"	)	,
(	"1001111011"	)	,
(	"1001111110"	)	,
(	"1010000001"	)	,
(	"1010000100"	)	,
(	"1010000111"	)	,
(	"1010001010"	)	,
(	"1010001101"	)	,
(	"1010010000"	)	,
(	"1010010011"	)	,
(	"1010010110"	)	,
(	"1010011001"	)	,
(	"1010011100"	)	,
(	"1010011111"	)	,
(	"1010100010"	)	,
(	"1010100101"	)	,
(	"1010101000"	)	,
(	"1010101011"	)	,
(	"1010101110"	)	,
(	"1010110001"	)	,
(	"1010110011"	)	,
(	"1010110110"	)	,
(	"1010111001"	)	,
(	"1010111100"	)	,
(	"1010111111"	)	,
(	"1011000010"	)	,
(	"1011000101"	)	,
(	"1011001000"	)	,
(	"1011001011"	)	,
(	"1011001110"	)	,
(	"1011010000"	)	,
(	"1011010011"	)	,
(	"1011010110"	)	,
(	"1011011001"	)	,
(	"1011011100"	)	,
(	"1011011111"	)	,
(	"1011100001"	)	,
(	"1011100100"	)	,
(	"1011100111"	)	,
(	"1011101010"	)	,
(	"1011101101"	)	,
(	"1011101111"	)	,
(	"1011110010"	)	,
(	"1011110101"	)	,
(	"1011111000"	)	,
(	"1011111010"	)	,
(	"1011111101"	)	,
(	"1100000000"	)	,
(	"1100000011"	)	,
(	"1100000101"	)	,
(	"1100001000"	)	,
(	"1100001011"	)	,
(	"1100001101"	)	,
(	"1100010000"	)	,
(	"1100010011"	)	,
(	"1100010101"	)	,
(	"1100011000"	)	,
(	"1100011010"	)	,
(	"1100011101"	)	,
(	"1100100000"	)	,
(	"1100100010"	)	,
(	"1100100101"	)	,
(	"1100100111"	)	,
(	"1100101010"	)	,
(	"1100101100"	)	,
(	"1100101111"	)	,
(	"1100110001"	)	,
(	"1100110100"	)	,
(	"1100110110"	)	,
(	"1100111001"	)	,
(	"1100111011"	)	,
(	"1100111110"	)	,
(	"1101000000"	)	,
(	"1101000011"	)	,
(	"1101000101"	)	,
(	"1101000111"	)	,
(	"1101001010"	)	,
(	"1101001100"	)	,
(	"1101001111"	)	,
(	"1101010001"	)	,
(	"1101010011"	)	,
(	"1101010110"	)	,
(	"1101011000"	)	,
(	"1101011010"	)	,
(	"1101011101"	)	,
(	"1101011111"	)	,
(	"1101100001"	)	,
(	"1101100011"	)	,
(	"1101100110"	)	,
(	"1101101000"	)	,
(	"1101101010"	)	,
(	"1101101100"	)	,
(	"1101101110"	)	,
(	"1101110001"	)	,
(	"1101110011"	)	,
(	"1101110101"	)	,
(	"1101110111"	)	,
(	"1101111001"	)	,
(	"1101111011"	)	,
(	"1101111101"	)	,
(	"1101111111"	)	,
(	"1110000001"	)	,
(	"1110000011"	)	,
(	"1110000110"	)	,
(	"1110001000"	)	,
(	"1110001010"	)	,
(	"1110001011"	)	,
(	"1110001101"	)	,
(	"1110001111"	)	,
(	"1110010001"	)	,
(	"1110010011"	)	,
(	"1110010101"	)	,
(	"1110010111"	)	,
(	"1110011001"	)	,
(	"1110011011"	)	,
(	"1110011101"	)	,
(	"1110011110"	)	,
(	"1110100000"	)	,
(	"1110100010"	)	,
(	"1110100100"	)	,
(	"1110100110"	)	,
(	"1110100111"	)	,
(	"1110101001"	)	,
(	"1110101011"	)	,
(	"1110101101"	)	,
(	"1110101110"	)	,
(	"1110110000"	)	,
(	"1110110010"	)	,
(	"1110110011"	)	,
(	"1110110101"	)	,
(	"1110110110"	)	,
(	"1110111000"	)	,
(	"1110111010"	)	,
(	"1110111011"	)	,
(	"1110111101"	)	,
(	"1110111110"	)	,
(	"1111000000"	)	,
(	"1111000001"	)	,
(	"1111000011"	)	,
(	"1111000100"	)	,
(	"1111000110"	)	,
(	"1111000111"	)	,
(	"1111001000"	)	,
(	"1111001010"	)	,
(	"1111001011"	)	,
(	"1111001100"	)	,
(	"1111001110"	)	,
(	"1111001111"	)	,
(	"1111010000"	)	,
(	"1111010010"	)	,
(	"1111010011"	)	,
(	"1111010100"	)	,
(	"1111010101"	)	,
(	"1111010111"	)	,
(	"1111011000"	)	,
(	"1111011001"	)	,
(	"1111011010"	)	,
(	"1111011011"	)	,
(	"1111011100"	)	,
(	"1111011101"	)	,
(	"1111011111"	)	,
(	"1111100000"	)	,
(	"1111100001"	)	,
(	"1111100010"	)	,
(	"1111100011"	)	,
(	"1111100100"	)	,
(	"1111100101"	)	,
(	"1111100110"	)	,
(	"1111100111"	)	,
(	"1111100111"	)	,
(	"1111101000"	)	,
(	"1111101001"	)	,
(	"1111101010"	)	,
(	"1111101011"	)	,
(	"1111101100"	)	,
(	"1111101101"	)	,
(	"1111101101"	)	,
(	"1111101110"	)	,
(	"1111101111"	)	,
(	"1111110000"	)	,
(	"1111110000"	)	,
(	"1111110001"	)	,
(	"1111110010"	)	,
(	"1111110010"	)	,
(	"1111110011"	)	,
(	"1111110100"	)	,
(	"1111110100"	)	,
(	"1111110101"	)	,
(	"1111110101"	)	,
(	"1111110110"	)	,
(	"1111110111"	)	,
(	"1111110111"	)	,
(	"1111110111"	)	,
(	"1111111000"	)	,
(	"1111111000"	)	,
(	"1111111001"	)	,
(	"1111111001"	)	,
(	"1111111010"	)	,
(	"1111111010"	)	,
(	"1111111010"	)	,
(	"1111111011"	)	,
(	"1111111011"	)	,
(	"1111111011"	)	,
(	"1111111100"	)	,
(	"1111111100"	)	,
(	"1111111100"	)	,
(	"1111111100"	)	,
(	"1111111101"	)	,
(	"1111111101"	)	,
(	"1111111101"	)	,
(	"1111111101"	)	,
(	"1111111101"	)	,
(	"1111111101"	)	,
(	"1111111101"	)	,
(	"1111111101"	)	,
(	"1111111101"	)	,
(	"1111111101"	)	,
(	"1111111110"	)	,
(	"1111111101"	)	,
(	"1111111101"	)	,
(	"1111111101"	)	,
(	"1111111101"	)	,
(	"1111111101"	)	,
(	"1111111101"	)	,
(	"1111111101"	)	,
(	"1111111101"	)	,
(	"1111111101"	)	,
(	"1111111101"	)	,
(	"1111111100"	)	,
(	"1111111100"	)	,
(	"1111111100"	)	,
(	"1111111100"	)	,
(	"1111111011"	)	,
(	"1111111011"	)	,
(	"1111111011"	)	,
(	"1111111010"	)	,
(	"1111111010"	)	,
(	"1111111010"	)	,
(	"1111111001"	)	,
(	"1111111001"	)	,
(	"1111111000"	)	,
(	"1111111000"	)	,
(	"1111110111"	)	,
(	"1111110111"	)	,
(	"1111110111"	)	,
(	"1111110110"	)	,
(	"1111110101"	)	,
(	"1111110101"	)	,
(	"1111110100"	)	,
(	"1111110100"	)	,
(	"1111110011"	)	,
(	"1111110010"	)	,
(	"1111110010"	)	,
(	"1111110001"	)	,
(	"1111110000"	)	,
(	"1111110000"	)	,
(	"1111101111"	)	,
(	"1111101110"	)	,
(	"1111101101"	)	,
(	"1111101101"	)	,
(	"1111101100"	)	,
(	"1111101011"	)	,
(	"1111101010"	)	,
(	"1111101001"	)	,
(	"1111101000"	)	,
(	"1111100111"	)	,
(	"1111100111"	)	,
(	"1111100110"	)	,
(	"1111100101"	)	,
(	"1111100100"	)	,
(	"1111100011"	)	,
(	"1111100010"	)	,
(	"1111100001"	)	,
(	"1111100000"	)	,
(	"1111011111"	)	,
(	"1111011101"	)	,
(	"1111011100"	)	,
(	"1111011011"	)	,
(	"1111011010"	)	,
(	"1111011001"	)	,
(	"1111011000"	)	,
(	"1111010111"	)	,
(	"1111010101"	)	,
(	"1111010100"	)	,
(	"1111010011"	)	,
(	"1111010010"	)	,
(	"1111010000"	)	,
(	"1111001111"	)	,
(	"1111001110"	)	,
(	"1111001100"	)	,
(	"1111001011"	)	,
(	"1111001010"	)	,
(	"1111001000"	)	,
(	"1111000111"	)	,
(	"1111000110"	)	,
(	"1111000100"	)	,
(	"1111000011"	)	,
(	"1111000001"	)	,
(	"1111000000"	)	,
(	"1110111110"	)	,
(	"1110111101"	)	,
(	"1110111011"	)	,
(	"1110111010"	)	,
(	"1110111000"	)	,
(	"1110110110"	)	,
(	"1110110101"	)	,
(	"1110110011"	)	,
(	"1110110010"	)	,
(	"1110110000"	)	,
(	"1110101110"	)	,
(	"1110101101"	)	,
(	"1110101011"	)	,
(	"1110101001"	)	,
(	"1110100111"	)	,
(	"1110100110"	)	,
(	"1110100100"	)	,
(	"1110100010"	)	,
(	"1110100000"	)	,
(	"1110011110"	)	,
(	"1110011101"	)	,
(	"1110011011"	)	,
(	"1110011001"	)	,
(	"1110010111"	)	,
(	"1110010101"	)	,
(	"1110010011"	)	,
(	"1110010001"	)	,
(	"1110001111"	)	,
(	"1110001101"	)	,
(	"1110001011"	)	,
(	"1110001010"	)	,
(	"1110001000"	)	,
(	"1110000110"	)	,
(	"1110000011"	)	,
(	"1110000001"	)	,
(	"1101111111"	)	,
(	"1101111101"	)	,
(	"1101111011"	)	,
(	"1101111001"	)	,
(	"1101110111"	)	,
(	"1101110101"	)	,
(	"1101110011"	)	,
(	"1101110001"	)	,
(	"1101101110"	)	,
(	"1101101100"	)	,
(	"1101101010"	)	,
(	"1101101000"	)	,
(	"1101100110"	)	,
(	"1101100011"	)	,
(	"1101100001"	)	,
(	"1101011111"	)	,
(	"1101011101"	)	,
(	"1101011010"	)	,
(	"1101011000"	)	,
(	"1101010110"	)	,
(	"1101010011"	)	,
(	"1101010001"	)	,
(	"1101001111"	)	,
(	"1101001100"	)	,
(	"1101001010"	)	,
(	"1101000111"	)	,
(	"1101000101"	)	,
(	"1101000011"	)	,
(	"1101000000"	)	,
(	"1100111110"	)	,
(	"1100111011"	)	,
(	"1100111001"	)	,
(	"1100110110"	)	,
(	"1100110100"	)	,
(	"1100110001"	)	,
(	"1100101111"	)	,
(	"1100101100"	)	,
(	"1100101010"	)	,
(	"1100100111"	)	,
(	"1100100101"	)	,
(	"1100100010"	)	,
(	"1100100000"	)	,
(	"1100011101"	)	,
(	"1100011010"	)	,
(	"1100011000"	)	,
(	"1100010101"	)	,
(	"1100010011"	)	,
(	"1100010000"	)	,
(	"1100001101"	)	,
(	"1100001011"	)	,
(	"1100001000"	)	,
(	"1100000101"	)	,
(	"1100000011"	)	,
(	"1100000000"	)	,
(	"1011111101"	)	,
(	"1011111010"	)	,
(	"1011111000"	)	,
(	"1011110101"	)	,
(	"1011110010"	)	,
(	"1011101111"	)	,
(	"1011101101"	)	,
(	"1011101010"	)	,
(	"1011100111"	)	,
(	"1011100100"	)	,
(	"1011100001"	)	,
(	"1011011111"	)	,
(	"1011011100"	)	,
(	"1011011001"	)	,
(	"1011010110"	)	,
(	"1011010011"	)	,
(	"1011010000"	)	,
(	"1011001110"	)	,
(	"1011001011"	)	,
(	"1011001000"	)	,
(	"1011000101"	)	,
(	"1011000010"	)	,
(	"1010111111"	)	,
(	"1010111100"	)	,
(	"1010111001"	)	,
(	"1010110110"	)	,
(	"1010110011"	)	,
(	"1010110001"	)	,
(	"1010101110"	)	,
(	"1010101011"	)	,
(	"1010101000"	)	,
(	"1010100101"	)	,
(	"1010100010"	)	,
(	"1010011111"	)	,
(	"1010011100"	)	,
(	"1010011001"	)	,
(	"1010010110"	)	,
(	"1010010011"	)	,
(	"1010010000"	)	,
(	"1010001101"	)	,
(	"1010001010"	)	,
(	"1010000111"	)	,
(	"1010000100"	)	,
(	"1010000001"	)	,
(	"1001111110"	)	,
(	"1001111011"	)	,
(	"1001111000"	)	,
(	"1001110101"	)	,
(	"1001110010"	)	,
(	"1001101110"	)	,
(	"1001101011"	)	,
(	"1001101000"	)	,
(	"1001100101"	)	,
(	"1001100010"	)	,
(	"1001011111"	)	,
(	"1001011100"	)	,
(	"1001011001"	)	,
(	"1001010110"	)	,
(	"1001010011"	)	,
(	"1001010000"	)	,
(	"1001001101"	)	,
(	"1001001001"	)	,
(	"1001000110"	)	,
(	"1001000011"	)	,
(	"1001000000"	)	,
(	"1000111101"	)	,
(	"1000111010"	)	,
(	"1000110111"	)	,
(	"1000110100"	)	,
(	"1000110001"	)	,
(	"1000101101"	)	,
(	"1000101010"	)	,
(	"1000100111"	)	,
(	"1000100100"	)	,
(	"1000100001"	)	,
(	"1000011110"	)	,
(	"1000011011"	)	,
(	"1000011000"	)	,
(	"1000010100"	)	,
(	"1000010001"	)	,
(	"1000001110"	)	,
(	"1000001011"	)	,
(	"1000001000"	)	,
(	"1000000101"	)	,
(	"1000000010"	)	,
(	"0111111111"	)	,
(	"0111111011"	)	,
(	"0111111000"	)	,
(	"0111110101"	)	,
(	"0111110010"	)	,
(	"0111101111"	)	,
(	"0111101100"	)	,
(	"0111101001"	)	,
(	"0111100101"	)	,
(	"0111100010"	)	,
(	"0111011111"	)	,
(	"0111011100"	)	,
(	"0111011001"	)	,
(	"0111010110"	)	,
(	"0111010011"	)	,
(	"0111010000"	)	,
(	"0111001100"	)	,
(	"0111001001"	)	,
(	"0111000110"	)	,
(	"0111000011"	)	,
(	"0111000000"	)	,
(	"0110111101"	)	,
(	"0110111010"	)	,
(	"0110110111"	)	,
(	"0110110100"	)	,
(	"0110110000"	)	,
(	"0110101101"	)	,
(	"0110101010"	)	,
(	"0110100111"	)	,
(	"0110100100"	)	,
(	"0110100001"	)	,
(	"0110011110"	)	,
(	"0110011011"	)	,
(	"0110011000"	)	,
(	"0110010101"	)	,
(	"0110010010"	)	,
(	"0110001111"	)	,
(	"0110001011"	)	,
(	"0110001000"	)	,
(	"0110000101"	)	,
(	"0110000010"	)	,
(	"0101111111"	)	,
(	"0101111100"	)	,
(	"0101111001"	)	,
(	"0101110110"	)	,
(	"0101110011"	)	,
(	"0101110000"	)	,
(	"0101101101"	)	,
(	"0101101010"	)	,
(	"0101100111"	)	,
(	"0101100100"	)	,
(	"0101100001"	)	,
(	"0101011110"	)	,
(	"0101011011"	)	,
(	"0101011000"	)	,
(	"0101010101"	)	,
(	"0101010010"	)	,
(	"0101001111"	)	,
(	"0101001100"	)	,
(	"0101001010"	)	,
(	"0101000111"	)	,
(	"0101000100"	)	,
(	"0101000001"	)	,
(	"0100111110"	)	,
(	"0100111011"	)	,
(	"0100111000"	)	,
(	"0100110101"	)	,
(	"0100110010"	)	,
(	"0100101111"	)	,
(	"0100101101"	)	,
(	"0100101010"	)	,
(	"0100100111"	)	,
(	"0100100100"	)	,
(	"0100100001"	)	,
(	"0100011110"	)	,
(	"0100011100"	)	,
(	"0100011001"	)	,
(	"0100010110"	)	,
(	"0100010011"	)	,
(	"0100010000"	)	,
(	"0100001110"	)	,
(	"0100001011"	)	,
(	"0100001000"	)	,
(	"0100000101"	)	,
(	"0100000011"	)	,
(	"0100000000"	)	,
(	"0011111101"	)	,
(	"0011111010"	)	,
(	"0011111000"	)	,
(	"0011110101"	)	,
(	"0011110010"	)	,
(	"0011110000"	)	,
(	"0011101101"	)	,
(	"0011101010"	)	,
(	"0011101000"	)	,
(	"0011100101"	)	,
(	"0011100011"	)	,
(	"0011100000"	)	,
(	"0011011101"	)	,
(	"0011011011"	)	,
(	"0011011000"	)	,
(	"0011010110"	)	,
(	"0011010011"	)	,
(	"0011010001"	)	,
(	"0011001110"	)	,
(	"0011001100"	)	,
(	"0011001001"	)	,
(	"0011000111"	)	,
(	"0011000100"	)	,
(	"0011000010"	)	,
(	"0010111111"	)	,
(	"0010111101"	)	,
(	"0010111010"	)	,
(	"0010111000"	)	,
(	"0010110110"	)	,
(	"0010110011"	)	,
(	"0010110001"	)	,
(	"0010101110"	)	,
(	"0010101100"	)	,
(	"0010101010"	)	,
(	"0010100111"	)	,
(	"0010100101"	)	,
(	"0010100011"	)	,
(	"0010100000"	)	,
(	"0010011110"	)	,
(	"0010011100"	)	,
(	"0010011010"	)	,
(	"0010010111"	)	,
(	"0010010101"	)	,
(	"0010010011"	)	,
(	"0010010001"	)	,
(	"0010001111"	)	,
(	"0010001100"	)	,
(	"0010001010"	)	,
(	"0010001000"	)	,
(	"0010000110"	)	,
(	"0010000100"	)	,
(	"0010000010"	)	,
(	"0010000000"	)	,
(	"0001111110"	)	,
(	"0001111100"	)	,
(	"0001111010"	)	,
(	"0001110111"	)	,
(	"0001110101"	)	,
(	"0001110011"	)	,
(	"0001110010"	)	,
(	"0001110000"	)	,
(	"0001101110"	)	,
(	"0001101100"	)	,
(	"0001101010"	)	,
(	"0001101000"	)	,
(	"0001100110"	)	,
(	"0001100100"	)	,
(	"0001100010"	)	,
(	"0001100000"	)	,
(	"0001011111"	)	,
(	"0001011101"	)	,
(	"0001011011"	)	,
(	"0001011001"	)	,
(	"0001010111"	)	,
(	"0001010110"	)	,
(	"0001010100"	)	,
(	"0001010010"	)	,
(	"0001010000"	)	,
(	"0001001111"	)	,
(	"0001001101"	)	,
(	"0001001011"	)	,
(	"0001001010"	)	,
(	"0001001000"	)	,
(	"0001000111"	)	,
(	"0001000101"	)	,
(	"0001000011"	)	,
(	"0001000010"	)	,
(	"0001000000"	)	,
(	"0000111111"	)	,
(	"0000111101"	)	,
(	"0000111100"	)	,
(	"0000111010"	)	,
(	"0000111001"	)	,
(	"0000110111"	)	,
(	"0000110110"	)	,
(	"0000110101"	)	,
(	"0000110011"	)	,
(	"0000110010"	)	,
(	"0000110001"	)	,
(	"0000101111"	)	,
(	"0000101110"	)	,
(	"0000101101"	)	,
(	"0000101011"	)	,
(	"0000101010"	)	,
(	"0000101001"	)	,
(	"0000101000"	)	,
(	"0000100110"	)	,
(	"0000100101"	)	,
(	"0000100100"	)	,
(	"0000100011"	)	,
(	"0000100010"	)	,
(	"0000100001"	)	,
(	"0000100000"	)	,
(	"0000011110"	)	,
(	"0000011101"	)	,
(	"0000011100"	)	,
(	"0000011011"	)	,
(	"0000011010"	)	,
(	"0000011001"	)	,
(	"0000011000"	)	,
(	"0000010111"	)	,
(	"0000010110"	)	,
(	"0000010110"	)	,
(	"0000010101"	)	,
(	"0000010100"	)	,
(	"0000010011"	)	,
(	"0000010010"	)	,
(	"0000010001"	)	,
(	"0000010000"	)	,
(	"0000010000"	)	,
(	"0000001111"	)	,
(	"0000001110"	)	,
(	"0000001101"	)	,
(	"0000001101"	)	,
(	"0000001100"	)	,
(	"0000001011"	)	,
(	"0000001011"	)	,
(	"0000001010"	)	,
(	"0000001001"	)	,
(	"0000001001"	)	,
(	"0000001000"	)	,
(	"0000001000"	)	,
(	"0000000111"	)	,
(	"0000000110"	)	,
(	"0000000110"	)	,
(	"0000000110"	)	,
(	"0000000101"	)	,
(	"0000000101"	)	,
(	"0000000100"	)	,
(	"0000000100"	)	,
(	"0000000011"	)	,
(	"0000000011"	)	,
(	"0000000011"	)	,
(	"0000000010"	)	,
(	"0000000010"	)	,
(	"0000000010"	)	,
(	"0000000001"	)	,
(	"0000000001"	)	,
(	"0000000001"	)	,
(	"0000000001"	)	,
(	"0000000000"	)	,
(	"0000000000"	)	,
(	"0000000000"	)	,
(	"0000000000"	)	,
(	"0000000000"	)	,
(	"0000000000"	)	,
(	"0000000000"	)	,
(	"0000000000"	)	,
(	"0000000000"	)	,
(	"0000000000"	)	,
(	"0000000000"	)	,
(	"0000000000"	)	,
(	"0000000000"	)	,
(	"0000000000"	)	,
(	"0000000000"	)	,
(	"0000000000"	)	,
(	"0000000000"	)	,
(	"0000000000"	)	,
(	"0000000000"	)	,
(	"0000000000"	)	,
(	"0000000000"	)	,
(	"0000000001"	)	,
(	"0000000001"	)	,
(	"0000000001"	)	,
(	"0000000001"	)	,
(	"0000000010"	)	,
(	"0000000010"	)	,
(	"0000000010"	)	,
(	"0000000011"	)	,
(	"0000000011"	)	,
(	"0000000011"	)	,
(	"0000000100"	)	,
(	"0000000100"	)	,
(	"0000000101"	)	,
(	"0000000101"	)	,
(	"0000000110"	)	,
(	"0000000110"	)	,
(	"0000000110"	)	,
(	"0000000111"	)	,
(	"0000001000"	)	,
(	"0000001000"	)	,
(	"0000001001"	)	,
(	"0000001001"	)	,
(	"0000001010"	)	,
(	"0000001011"	)	,
(	"0000001011"	)	,
(	"0000001100"	)	,
(	"0000001101"	)	,
(	"0000001101"	)	,
(	"0000001110"	)	,
(	"0000001111"	)	,
(	"0000010000"	)	,
(	"0000010000"	)	,
(	"0000010001"	)	,
(	"0000010010"	)	,
(	"0000010011"	)	,
(	"0000010100"	)	,
(	"0000010101"	)	,
(	"0000010110"	)	,
(	"0000010110"	)	,
(	"0000010111"	)	,
(	"0000011000"	)	,
(	"0000011001"	)	,
(	"0000011010"	)	,
(	"0000011011"	)	,
(	"0000011100"	)	,
(	"0000011101"	)	,
(	"0000011110"	)	,
(	"0000100000"	)	,
(	"0000100001"	)	,
(	"0000100010"	)	,
(	"0000100011"	)	,
(	"0000100100"	)	,
(	"0000100101"	)	,
(	"0000100110"	)	,
(	"0000101000"	)	,
(	"0000101001"	)	,
(	"0000101010"	)	,
(	"0000101011"	)	,
(	"0000101101"	)	,
(	"0000101110"	)	,
(	"0000101111"	)	,
(	"0000110001"	)	,
(	"0000110010"	)	,
(	"0000110011"	)	,
(	"0000110101"	)	,
(	"0000110110"	)	,
(	"0000110111"	)	,
(	"0000111001"	)	,
(	"0000111010"	)	,
(	"0000111100"	)	,
(	"0000111101"	)	,
(	"0000111111"	)	,
(	"0001000000"	)	,
(	"0001000010"	)	,
(	"0001000011"	)	,
(	"0001000101"	)	,
(	"0001000111"	)	,
(	"0001001000"	)	,
(	"0001001010"	)	,
(	"0001001011"	)	,
(	"0001001101"	)	,
(	"0001001111"	)	,
(	"0001010000"	)	,
(	"0001010010"	)	,
(	"0001010100"	)	,
(	"0001010110"	)	,
(	"0001010111"	)	,
(	"0001011001"	)	,
(	"0001011011"	)	,
(	"0001011101"	)	,
(	"0001011111"	)	,
(	"0001100000"	)	,
(	"0001100010"	)	,
(	"0001100100"	)	,
(	"0001100110"	)	,
(	"0001101000"	)	,
(	"0001101010"	)	,
(	"0001101100"	)	,
(	"0001101110"	)	,
(	"0001110000"	)	,
(	"0001110010"	)	,
(	"0001110011"	)	,
(	"0001110101"	)	,
(	"0001110111"	)	,
(	"0001111010"	)	,
(	"0001111100"	)	,
(	"0001111110"	)	,
(	"0010000000"	)	,
(	"0010000010"	)	,
(	"0010000100"	)	,
(	"0010000110"	)	,
(	"0010001000"	)	,
(	"0010001010"	)	,
(	"0010001100"	)	,
(	"0010001111"	)	,
(	"0010010001"	)	,
(	"0010010011"	)	,
(	"0010010101"	)	,
(	"0010010111"	)	,
(	"0010011010"	)	,
(	"0010011100"	)	,
(	"0010011110"	)	,
(	"0010100000"	)	,
(	"0010100011"	)	,
(	"0010100101"	)	,
(	"0010100111"	)	,
(	"0010101010"	)	,
(	"0010101100"	)	,
(	"0010101110"	)	,
(	"0010110001"	)	,
(	"0010110011"	)	,
(	"0010110110"	)	,
(	"0010111000"	)	,
(	"0010111010"	)	,
(	"0010111101"	)	,
(	"0010111111"	)	,
(	"0011000010"	)	,
(	"0011000100"	)	,
(	"0011000111"	)	,
(	"0011001001"	)	,
(	"0011001100"	)	,
(	"0011001110"	)	,
(	"0011010001"	)	,
(	"0011010011"	)	,
(	"0011010110"	)	,
(	"0011011000"	)	,
(	"0011011011"	)	,
(	"0011011101"	)	,
(	"0011100000"	)	,
(	"0011100011"	)	,
(	"0011100101"	)	,
(	"0011101000"	)	,
(	"0011101010"	)	,
(	"0011101101"	)	,
(	"0011110000"	)	,
(	"0011110010"	)	,
(	"0011110101"	)	,
(	"0011111000"	)	,
(	"0011111010"	)	,
(	"0011111101"	)	,
(	"0100000000"	)	,
(	"0100000011"	)	,
(	"0100000101"	)	,
(	"0100001000"	)	,
(	"0100001011"	)	,
(	"0100001110"	)	,
(	"0100010000"	)	,
(	"0100010011"	)	,
(	"0100010110"	)	,
(	"0100011001"	)	,
(	"0100011100"	)	,
(	"0100011110"	)	,
(	"0100100001"	)	,
(	"0100100100"	)	,
(	"0100100111"	)	,
(	"0100101010"	)	,
(	"0100101101"	)	,
(	"0100101111"	)	,
(	"0100110010"	)	,
(	"0100110101"	)	,
(	"0100111000"	)	,
(	"0100111011"	)	,
(	"0100111110"	)	,
(	"0101000001"	)	,
(	"0101000100"	)	,
(	"0101000111"	)	,
(	"0101001010"	)	,
(	"0101001100"	)	,
(	"0101001111"	)	,
(	"0101010010"	)	,
(	"0101010101"	)	,
(	"0101011000"	)	,
(	"0101011011"	)	,
(	"0101011110"	)	,
(	"0101100001"	)	,
(	"0101100100"	)	,
(	"0101100111"	)	,
(	"0101101010"	)	,
(	"0101101101"	)	,
(	"0101110000"	)	,
(	"0101110011"	)	,
(	"0101110110"	)	,
(	"0101111001"	)	,
(	"0101111100"	)	,
(	"0101111111"	)	,
(	"0110000010"	)	,
(	"0110000101"	)	,
(	"0110001000"	)	,
(	"0110001011"	)	,
(	"0110001111"	)	,
(	"0110010010"	)	,
(	"0110010101"	)	,
(	"0110011000"	)	,
(	"0110011011"	)	,
(	"0110011110"	)	,
(	"0110100001"	)	,
(	"0110100100"	)	,
(	"0110100111"	)	,
(	"0110101010"	)	,
(	"0110101101"	)	,
(	"0110110000"	)	,
(	"0110110100"	)	,
(	"0110110111"	)	,
(	"0110111010"	)	,
(	"0110111101"	)	,
(	"0111000000"	)	,
(	"0111000011"	)	,
(	"0111000110"	)	,
(	"0111001001"	)	,
(	"0111001100"	)	,
(	"0111010000"	)	,
(	"0111010011"	)	,
(	"0111010110"	)	,
(	"0111011001"	)	,
(	"0111011100"	)	,
(	"0111011111"	)	,
(	"0111100010"	)	,
(	"0111100101"	)	,
(	"0111101001"	)	,
(	"0111101100"	)	,
(	"0111101111"	)	,
(	"0111110010"	)	,
(	"0111110101"	)	,
(	"0111111000"	)	,
(	"0111111011"	)
);


begin
	
	yeet : process(index)
	begin
		if(index < 0) then
			duty_cycle <= "0000000000";
		elsif (index > 4095) then
			duty_cycle <= "0000000000";
		else
			duty_cycle <= Sinevalues(index);
		end if;
	end process;
--	duty_cycle <= std_logic_vector(to_unsigned(sawtooth(to_integer(unsigned(index))),duty_cycle'length));

end behavior;
