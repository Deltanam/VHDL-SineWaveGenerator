 
-- In this example, we're going to map voltage to distance, using a linear 
-- approximation, according to the Sharp GP2Y0A41SK0F datasheet page 4, or 
-- Lab 3 handout page 5. 
-- 
-- The relevant points we will select are:
-- 2.750 V is  4.00 cm (or 2750 mV and  40.0 mm)
-- 0.400 V is 33.00 cm (or  400 mV and 330.0 mm)
-- 
-- Mapping to the scales in our system
-- 2750 (mV) should map to  400 (10^-4 m)
--  400 (mV) should map to 3300 (10^-4 m)
-- and developing a linear equation, we find:
--
-- Distance = -2900/2350 * Voltage + 3793.617
-- Note this code implements linear function, you must map to the 
-- NON-linear relationship in the datasheet. This code is only provided 
-- for reference to help get you started.

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY BuzzAmp_Lookup IS
   PORT(
      clk            :  IN    STD_LOGIC;                                
      reset          :  IN    STD_LOGIC;                                
      index      	 :  IN    integer;                           
      Amplitude     :  OUT   integer
		);
END BuzzAmp_Lookup;

ARCHITECTURE behavior OF BuzzAmp_Lookup IS

type array_1d is array (0 to 4095) of integer;

constant BuzzAmps : array_1d := (				
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4093),
(4092),
(4090),
(4088),
(4087),
(4085),
(4083),
(4082),
(4080),
(4078),
(4077),
(4075),
(4073),
(4072),
(4070),
(4069),
(4067),
(4065),
(4064),
(4062),
(4060),
(4059),
(4057),
(4055),
(4054),
(4052),
(4050),
(4049),
(4047),
(4045),
(4044),
(4042),
(4040),
(4039),
(4037),
(4035),
(4034),
(4032),
(4030),
(4029),
(4027),
(4025),
(4024),
(4022),
(4021),
(4019),
(4017),
(4016),
(4014),
(4012),
(4011),
(4009),
(4007),
(4006),
(4004),
(4002),
(4001),
(3999),
(3997),
(3996),
(3994),
(3992),
(3991),
(3989),
(3987),
(3986),
(3984),
(3982),
(3981),
(3979),
(3977),
(3976),
(3974),
(3973),
(3971),
(3969),
(3968),
(3966),
(3964),
(3963),
(3961),
(3959),
(3958),
(3956),
(3954),
(3953),
(3951),
(3949),
(3948),
(3946),
(3944),
(3943),
(3941),
(3939),
(3938),
(3936),
(3934),
(3933),
(3931),
(3930),
(3928),
(3926),
(3925),
(3923),
(3921),
(3920),
(3918),
(3916),
(3915),
(3913),
(3911),
(3910),
(3908),
(3906),
(3905),
(3903),
(3901),
(3900),
(3898),
(3896),
(3895),
(3893),
(3891),
(3890),
(3888),
(3886),
(3885),
(3883),
(3882),
(3880),
(3878),
(3877),
(3875),
(3873),
(3872),
(3870),
(3868),
(3867),
(3865),
(3863),
(3862),
(3860),
(3858),
(3857),
(3855),
(3853),
(3852),
(3850),
(3848),
(3847),
(3845),
(3843),
(3842),
(3840),
(3838),
(3837),
(3835),
(3834),
(3832),
(3830),
(3829),
(3827),
(3825),
(3824),
(3822),
(3820),
(3819),
(3817),
(3815),
(3814),
(3812),
(3810),
(3809),
(3807),
(3805),
(3804),
(3802),
(3800),
(3799),
(3797),
(3795),
(3794),
(3792),
(3790),
(3789),
(3787),
(3786),
(3784),
(3782),
(3781),
(3779),
(3777),
(3776),
(3774),
(3772),
(3771),
(3769),
(3767),
(3766),
(3764),
(3762),
(3761),
(3759),
(3757),
(3756),
(3754),
(3752),
(3751),
(3749),
(3747),
(3746),
(3744),
(3742),
(3741),
(3739),
(3738),
(3736),
(3734),
(3733),
(3731),
(3729),
(3728),
(3726),
(3724),
(3723),
(3721),
(3719),
(3718),
(3716),
(3714),
(3713),
(3711),
(3709),
(3708),
(3706),
(3704),
(3703),
(3701),
(3699),
(3698),
(3696),
(3695),
(3693),
(3691),
(3690),
(3688),
(3686),
(3685),
(3683),
(3681),
(3680),
(3678),
(3676),
(3675),
(3673),
(3671),
(3670),
(3668),
(3666),
(3665),
(3663),
(3661),
(3660),
(3658),
(3656),
(3655),
(3653),
(3651),
(3650),
(3648),
(3647),
(3645),
(3643),
(3642),
(3640),
(3638),
(3637),
(3635),
(3633),
(3632),
(3630),
(3628),
(3627),
(3625),
(3623),
(3622),
(3620),
(3618),
(3617),
(3615),
(3613),
(3612),
(3610),
(3608),
(3607),
(3605),
(3603),
(3602),
(3600),
(3599),
(3597),
(3595),
(3594),
(3592),
(3590),
(3589),
(3587),
(3585),
(3584),
(3582),
(3580),
(3579),
(3577),
(3575),
(3574),
(3572),
(3570),
(3569),
(3567),
(3565),
(3564),
(3562),
(3560),
(3559),
(3557),
(3555),
(3554),
(3552),
(3551),
(3549),
(3547),
(3546),
(3544),
(3542),
(3541),
(3539),
(3537),
(3536),
(3534),
(3532),
(3531),
(3529),
(3527),
(3526),
(3524),
(3522),
(3521),
(3519),
(3517),
(3516),
(3514),
(3512),
(3511),
(3509),
(3507),
(3506),
(3504),
(3503),
(3501),
(3499),
(3498),
(3496),
(3494),
(3493),
(3491),
(3489),
(3488),
(3486),
(3484),
(3483),
(3481),
(3479),
(3478),
(3476),
(3474),
(3473),
(3471),
(3469),
(3468),
(3466),
(3464),
(3463),
(3461),
(3459),
(3458),
(3456),
(3455),
(3453),
(3451),
(3450),
(3448),
(3446),
(3445),
(3443),
(3441),
(3440),
(3438),
(3436),
(3435),
(3433),
(3431),
(3430),
(3428),
(3426),
(3425),
(3423),
(3421),
(3420),
(3418),
(3416),
(3415),
(3413),
(3412),
(3410),
(3408),
(3407),
(3405),
(3403),
(3402),
(3400),
(3398),
(3397),
(3395),
(3393),
(3392),
(3390),
(3388),
(3387),
(3385),
(3383),
(3382),
(3380),
(3378),
(3377),
(3375),
(3373),
(3372),
(3370),
(3368),
(3367),
(3365),
(3364),
(3362),
(3360),
(3359),
(3357),
(3355),
(3354),
(3352),
(3350),
(3349),
(3347),
(3345),
(3344),
(3342),
(3340),
(3339),
(3337),
(3335),
(3334),
(3332),
(3330),
(3329),
(3327),
(3325),
(3324),
(3322),
(3320),
(3319),
(3317),
(3316),
(3314),
(3312),
(3311),
(3309),
(3307),
(3306),
(3304),
(3302),
(3301),
(3299),
(3297),
(3296),
(3294),
(3292),
(3291),
(3289),
(3287),
(3286),
(3284),
(3282),
(3281),
(3279),
(3277),
(3276),
(3274),
(3272),
(3271),
(3269),
(3268),
(3266),
(3264),
(3263),
(3261),
(3259),
(3258),
(3256),
(3254),
(3253),
(3251),
(3249),
(3248),
(3246),
(3244),
(3243),
(3241),
(3239),
(3238),
(3236),
(3234),
(3233),
(3231),
(3229),
(3228),
(3226),
(3224),
(3223),
(3221),
(3220),
(3218),
(3216),
(3215),
(3213),
(3211),
(3210),
(3208),
(3206),
(3205),
(3203),
(3201),
(3200),
(3198),
(3196),
(3195),
(3193),
(3191),
(3190),
(3188),
(3186),
(3185),
(3183),
(3181),
(3180),
(3178),
(3177),
(3175),
(3173),
(3172),
(3170),
(3168),
(3167),
(3165),
(3163),
(3162),
(3160),
(3158),
(3157),
(3155),
(3153),
(3152),
(3150),
(3148),
(3147),
(3145),
(3143),
(3142),
(3140),
(3138),
(3137),
(3135),
(3133),
(3132),
(3130),
(3129),
(3127),
(3125),
(3124),
(3122),
(3120),
(3119),
(3117),
(3115),
(3114),
(3112),
(3110),
(3109),
(3107),
(3105),
(3104),
(3102),
(3100),
(3099),
(3097),
(3095),
(3094),
(3092),
(3090),
(3089),
(3087),
(3085),
(3084),
(3082),
(3081),
(3079),
(3077),
(3076),
(3074),
(3072),
(3071),
(3069),
(3067),
(3066),
(3064),
(3062),
(3061),
(3059),
(3057),
(3056),
(3054),
(3052),
(3051),
(3049),
(3047),
(3046),
(3044),
(3042),
(3041),
(3039),
(3037),
(3036),
(3034),
(3033),
(3031),
(3029),
(3028),
(3026),
(3024),
(3023),
(3021),
(3019),
(3018),
(3016),
(3014),
(3013),
(3011),
(3009),
(3008),
(3006),
(3004),
(3003),
(3001),
(2999),
(2998),
(2996),
(2994),
(2993),
(2991),
(2989),
(2988),
(2986),
(2985),
(2983),
(2981),
(2980),
(2978),
(2976),
(2975),
(2973),
(2971),
(2970),
(2968),
(2966),
(2965),
(2963),
(2961),
(2960),
(2958),
(2956),
(2955),
(2953),
(2951),
(2950),
(2948),
(2946),
(2945),
(2943),
(2942),
(2940),
(2938),
(2937),
(2935),
(2933),
(2932),
(2930),
(2928),
(2927),
(2925),
(2923),
(2922),
(2920),
(2918),
(2917),
(2915),
(2913),
(2912),
(2910),
(2908),
(2907),
(2905),
(2903),
(2902),
(2900),
(2898),
(2897),
(2895),
(2894),
(2892),
(2890),
(2889),
(2887),
(2885),
(2884),
(2882),
(2880),
(2879),
(2877),
(2875),
(2874),
(2872),
(2870),
(2869),
(2867),
(2865),
(2864),
(2862),
(2860),
(2859),
(2857),
(2855),
(2854),
(2852),
(2850),
(2849),
(2847),
(2846),
(2844),
(2842),
(2841),
(2839),
(2837),
(2836),
(2834),
(2832),
(2831),
(2829),
(2827),
(2826),
(2824),
(2822),
(2821),
(2819),
(2817),
(2816),
(2814),
(2812),
(2811),
(2809),
(2807),
(2806),
(2804),
(2802),
(2801),
(2799),
(2798),
(2796),
(2794),
(2793),
(2791),
(2789),
(2788),
(2786),
(2784),
(2783),
(2781),
(2779),
(2778),
(2776),
(2774),
(2773),
(2771),
(2769),
(2768),
(2766),
(2764),
(2763),
(2761),
(2759),
(2758),
(2756),
(2754),
(2753),
(2751),
(2750),
(2748),
(2746),
(2745),
(2743),
(2741),
(2740),
(2738),
(2736),
(2735),
(2733),
(2731),
(2730),
(2728),
(2726),
(2725),
(2723),
(2721),
(2720),
(2718),
(2716),
(2715),
(2713),
(2711),
(2710),
(2708),
(2706),
(2705),
(2703),
(2702),
(2700),
(2698),
(2697),
(2695),
(2693),
(2692),
(2690),
(2688),
(2687),
(2685),
(2683),
(2682),
(2680),
(2678),
(2677),
(2675),
(2673),
(2672),
(2670),
(2668),
(2667),
(2665),
(2663),
(2662),
(2660),
(2659),
(2657),
(2655),
(2654),
(2652),
(2650),
(2649),
(2647),
(2645),
(2644),
(2642),
(2640),
(2639),
(2637),
(2635),
(2634),
(2632),
(2630),
(2629),
(2627),
(2625),
(2624),
(2622),
(2620),
(2619),
(2617),
(2615),
(2614),
(2612),
(2611),
(2609),
(2607),
(2606),
(2604),
(2602),
(2601),
(2599),
(2597),
(2596),
(2594),
(2592),
(2591),
(2589),
(2587),
(2586),
(2584),
(2582),
(2581),
(2579),
(2577),
(2576),
(2574),
(2572),
(2571),
(2569),
(2567),
(2566),
(2564),
(2563),
(2561),
(2559),
(2558),
(2556),
(2554),
(2553),
(2551),
(2549),
(2548),
(2546),
(2544),
(2543),
(2541),
(2539),
(2538),
(2536),
(2534),
(2533),
(2531),
(2529),
(2528),
(2526),
(2524),
(2523),
(2521),
(2519),
(2518),
(2516),
(2515),
(2513),
(2511),
(2510),
(2508),
(2506),
(2505),
(2503),
(2501),
(2500),
(2498),
(2496),
(2495),
(2493),
(2491),
(2490),
(2488),
(2486),
(2485),
(2483),
(2481),
(2480),
(2478),
(2476),
(2475),
(2473),
(2471),
(2470),
(2468),
(2467),
(2465),
(2463),
(2462),
(2460),
(2458),
(2457),
(2455),
(2453),
(2452),
(2450),
(2448),
(2447),
(2445),
(2443),
(2442),
(2440),
(2438),
(2437),
(2435),
(2433),
(2432),
(2430),
(2428),
(2427),
(2425),
(2424),
(2422),
(2420),
(2419),
(2417),
(2415),
(2414),
(2412),
(2410),
(2409),
(2407),
(2405),
(2404),
(2402),
(2400),
(2399),
(2397),
(2395),
(2394),
(2392),
(2390),
(2389),
(2387),
(2385),
(2384),
(2382),
(2380),
(2379),
(2377),
(2376),
(2374),
(2372),
(2371),
(2369),
(2367),
(2366),
(2364),
(2362),
(2361),
(2359),
(2357),
(2356),
(2354),
(2352),
(2351),
(2349),
(2347),
(2346),
(2344),
(2342),
(2341),
(2339),
(2337),
(2336),
(2334),
(2332),
(2331),
(2329),
(2328),
(2326),
(2324),
(2323),
(2321),
(2319),
(2318),
(2316),
(2314),
(2313),
(2311),
(2309),
(2308),
(2306),
(2304),
(2303),
(2301),
(2299),
(2298),
(2296),
(2294),
(2293),
(2291),
(2289),
(2288),
(2286),
(2284),
(2283),
(2281),
(2280),
(2278),
(2276),
(2275),
(2273),
(2271),
(2270),
(2268),
(2266),
(2265),
(2263),
(2261),
(2260),
(2258),
(2256),
(2255),
(2253),
(2251),
(2250),
(2248),
(2246),
(2245),
(2243),
(2241),
(2240),
(2238),
(2236),
(2235),
(2233),
(2232),
(2230),
(2228),
(2227),
(2225),
(2223),
(2222),
(2220),
(2218),
(2217),
(2215),
(2213),
(2212),
(2210),
(2208),
(2207),
(2205),
(2203),
(2202),
(2200),
(2198),
(2197),
(2195),
(2193),
(2192),
(2190),
(2188),
(2187),
(2185),
(2184),
(2182),
(2180),
(2179),
(2177),
(2175),
(2174),
(2172),
(2170),
(2169),
(2167),
(2165),
(2164),
(2162),
(2160),
(2159),
(2157),
(2155),
(2154),
(2152),
(2150),
(2149),
(2147),
(2145),
(2144),
(2142),
(2141),
(2139),
(2137),
(2136),
(2134),
(2132),
(2131),
(2129),
(2127),
(2126),
(2124),
(2122),
(2121),
(2119),
(2117),
(2116),
(2114),
(2112),
(2111),
(2109),
(2107),
(2106),
(2104),
(2102),
(2101),
(2099),
(2097),
(2096),
(2094),
(2093),
(2091),
(2089),
(2088),
(2086),
(2084),
(2083),
(2081),
(2079),
(2078),
(2076),
(2074),
(2073),
(2071),
(2069),
(2068),
(2066),
(2064),
(2063),
(2061),
(2059),
(2058),
(2056),
(2054),
(2053),
(2051),
(2049),
(2048),
(2046),
(2045),
(2043),
(2041),
(2040),
(2038),
(2036),
(2035),
(2033),
(2031),
(2030),
(2028),
(2026),
(2025),
(2023),
(2021),
(2020),
(2018),
(2016),
(2015),
(2013),
(2011),
(2010),
(2008),
(2006),
(2005),
(2003),
(2001),
(2000),
(1998),
(1997),
(1995),
(1993),
(1992),
(1990),
(1988),
(1987),
(1985),
(1983),
(1982),
(1980),
(1978),
(1977),
(1975),
(1973),
(1972),
(1970),
(1968),
(1967),
(1965),
(1963),
(1962),
(1960),
(1958),
(1957),
(1955),
(1953),
(1952),
(1950),
(1949),
(1947),
(1945),
(1944),
(1942),
(1940),
(1939),
(1937),
(1935),
(1934),
(1932),
(1930),
(1929),
(1927),
(1925),
(1924),
(1922),
(1920),
(1919),
(1917),
(1915),
(1914),
(1912),
(1910),
(1909),
(1907),
(1906),
(1904),
(1902),
(1901),
(1899),
(1897),
(1896),
(1894),
(1892),
(1891),
(1889),
(1887),
(1886),
(1884),
(1882),
(1881),
(1879),
(1877),
(1876),
(1874),
(1872),
(1871),
(1869),
(1867),
(1866),
(1864),
(1862),
(1861),
(1859),
(1858),
(1856),
(1854),
(1853),
(1851),
(1849),
(1848),
(1846),
(1844),
(1843),
(1841),
(1839),
(1838),
(1836),
(1834),
(1833),
(1831),
(1829),
(1828),
(1826),
(1824),
(1823),
(1821),
(1819),
(1818),
(1816),
(1814),
(1813),
(1811),
(1810),
(1808),
(1806),
(1805),
(1803),
(1801),
(1800),
(1798),
(1796),
(1795),
(1793),
(1791),
(1790),
(1788),
(1786),
(1785),
(1783),
(1781),
(1780),
(1778),
(1776),
(1775),
(1773),
(1771),
(1770),
(1768),
(1766),
(1765),
(1763),
(1762),
(1760),
(1758),
(1757),
(1755),
(1753),
(1752),
(1750),
(1748),
(1747),
(1745),
(1743),
(1742),
(1740),
(1738),
(1737),
(1735),
(1733),
(1732),
(1730),
(1728),
(1727),
(1725),
(1723),
(1722),
(1720),
(1718),
(1717),
(1715),
(1714),
(1712),
(1710),
(1709),
(1707),
(1705),
(1704),
(1702),
(1700),
(1699),
(1697),
(1695),
(1694),
(1692),
(1690),
(1689),
(1687),
(1685),
(1684),
(1682),
(1680),
(1679),
(1677),
(1675),
(1674),
(1672),
(1670),
(1669),
(1667),
(1666),
(1664),
(1662),
(1661),
(1659),
(1657),
(1656),
(1654),
(1652),
(1651),
(1649),
(1647),
(1646),
(1644),
(1642),
(1641),
(1639),
(1637),
(1636),
(1634),
(1632),
(1631),
(1629),
(1627),
(1626),
(1624),
(1623),
(1621),
(1619),
(1618),
(1616),
(1614),
(1613),
(1611),
(1609),
(1608),
(1606),
(1604),
(1603),
(1601),
(1599),
(1598),
(1596),
(1594),
(1593),
(1591),
(1589),
(1588),
(1586),
(1584),
(1583),
(1581),
(1579),
(1578),
(1576),
(1575),
(1573),
(1571),
(1570),
(1568),
(1566),
(1565),
(1563),
(1561),
(1560),
(1558),
(1556),
(1555),
(1553),
(1551),
(1550),
(1548),
(1546),
(1545),
(1543),
(1541),
(1540),
(1538),
(1536),
(1535),
(1533),
(1531),
(1530),
(1528),
(1527),
(1525),
(1523),
(1522),
(1520),
(1518),
(1517),
(1515),
(1513),
(1512),
(1510),
(1508),
(1507),
(1505),
(1503),
(1502),
(1500),
(1498),
(1497),
(1495),
(1493),
(1492),
(1490),
(1488),
(1487),
(1485),
(1483),
(1482),
(1480),
(1479),
(1477),
(1475),
(1474),
(1472),
(1470),
(1469),
(1467),
(1465),
(1464),
(1462),
(1460),
(1459),
(1457),
(1455),
(1454),
(1452),
(1450),
(1449),
(1447),
(1445),
(1444),
(1442),
(1440),
(1439),
(1437),
(1435),
(1434),
(1432),
(1431),
(1429),
(1427),
(1426),
(1424),
(1422),
(1421),
(1419),
(1417),
(1416),
(1414),
(1412),
(1411),
(1409),
(1407),
(1406),
(1404),
(1402),
(1401),
(1399),
(1397),
(1396),
(1394),
(1392),
(1391),
(1389),
(1388),
(1386),
(1384),
(1383),
(1381),
(1379),
(1378),
(1376),
(1374),
(1373),
(1371),
(1369),
(1368),
(1366),
(1364),
(1363),
(1361),
(1359),
(1358),
(1356),
(1354),
(1353),
(1351),
(1349),
(1348),
(1346),
(1344),
(1343),
(1341),
(1340),
(1338),
(1336),
(1335),
(1333),
(1331),
(1330),
(1328),
(1326),
(1325),
(1323),
(1321),
(1320),
(1318),
(1316),
(1315),
(1313),
(1311),
(1310),
(1308),
(1306),
(1305),
(1303),
(1301),
(1300),
(1298),
(1296),
(1295),
(1293),
(1292),
(1290),
(1288),
(1287),
(1285),
(1283),
(1282),
(1280),
(1278),
(1277),
(1275),
(1273),
(1272),
(1270),
(1268),
(1267),
(1265),
(1263),
(1262),
(1260),
(1258),
(1257),
(1255),
(1253),
(1252),
(1250),
(1248),
(1247),
(1245),
(1244),
(1242),
(1240),
(1239),
(1237),
(1235),
(1234),
(1232),
(1230),
(1229),
(1227),
(1225),
(1224),
(1222),
(1220),
(1219),
(1217),
(1215),
(1214),
(1212),
(1210),
(1209),
(1207),
(1205),
(1204),
(1202),
(1200),
(1199),
(1197),
(1196),
(1194),
(1192),
(1191),
(1189),
(1187),
(1186),
(1184),
(1182),
(1181),
(1179),
(1177),
(1176),
(1174),
(1172),
(1171),
(1169),
(1167),
(1166),
(1164),
(1162),
(1161),
(1159),
(1157),
(1156),
(1154),
(1152),
(1151),
(1149),
(1148),
(1146),
(1144),
(1143),
(1141),
(1139),
(1138),
(1136),
(1134),
(1133),
(1131),
(1129),
(1128),
(1126),
(1124),
(1123),
(1121),
(1119),
(1118),
(1116),
(1114),
(1113),
(1111),
(1109),
(1108),
(1106),
(1105),
(1103),
(1101),
(1100),
(1098),
(1096),
(1095),
(1093),
(1091),
(1090),
(1088),
(1086),
(1085),
(1083),
(1081),
(1080),
(1078),
(1076),
(1075),
(1073),
(1071),
(1070),
(1068),
(1066),
(1065),
(1063),
(1061),
(1060),
(1058),
(1057),
(1055),
(1053),
(1052),
(1050),
(1048),
(1047),
(1045),
(1043),
(1042),
(1040),
(1038),
(1037),
(1035),
(1033),
(1032),
(1030),
(1028),
(1027),
(1025),
(1023),
(1022),
(1020),
(1018),
(1017),
(1015),
(1013),
(1012),
(1010),
(1009),
(1007),
(1005),
(1004),
(1002),
(1000),
(999),
(997),
(995),
(994),
(992),
(990),
(989),
(987),
(985),
(984),
(982),
(980),
(979),
(977),
(975),
(974),
(972),
(970),
(969),
(967),
(965),
(964),
(962),
(961),
(959),
(957),
(956),
(954),
(952),
(951),
(949),
(947),
(946),
(944),
(942),
(941),
(939),
(937),
(936),
(934),
(932),
(931),
(929),
(927),
(926),
(924),
(922),
(921),
(919),
(917),
(916),
(914),
(913),
(911),
(909),
(908),
(906),
(904),
(903),
(901),
(899),
(898),
(896),
(894),
(893),
(891),
(889),
(888),
(886),
(884),
(883),
(881),
(879),
(878),
(876),
(874),
(873),
(871),
(870),
(868),
(866),
(865),
(863),
(861),
(860),
(858),
(856),
(855),
(853),
(851),
(850),
(848),
(846),
(845),
(843),
(841),
(840),
(838),
(836),
(835),
(833),
(831),
(830),
(828),
(826),
(825),
(823),
(822),
(820),
(818),
(817),
(815),
(813),
(812),
(810),
(808),
(807),
(805),
(803),
(802),
(800),
(798),
(797),
(795),
(793),
(792),
(790),
(788),
(787),
(785),
(783),
(782),
(780),
(778),
(777),
(775),
(774),
(772),
(770),
(769),
(767),
(765),
(764),
(762),
(760),
(759),
(757),
(755),
(754),
(752),
(750),
(749),
(747),
(745),
(744),
(742),
(740),
(739),
(737),
(735),
(734),
(732),
(730),
(729),
(727),
(726),
(724),
(722),
(721),
(719),
(717),
(716),
(714),
(712),
(711),
(709),
(707),
(706),
(704),
(702),
(701),
(699),
(697),
(696),
(694),
(692),
(691),
(689),
(687),
(686),
(684),
(682),
(681),
(679),
(678),
(676),
(674),
(673),
(671),
(669),
(668),
(666),
(664),
(663),
(661),
(659),
(658),
(656),
(654),
(653),
(651),
(649),
(648),
(646),
(644),
(643),
(641),
(639),
(638),
(636),
(635),
(633),
(631),
(630),
(628),
(626),
(625),
(623),
(621),
(620),
(618),
(616),
(615),
(613),
(611),
(610),
(608),
(606),
(605),
(603),
(601),
(600),
(598),
(596),
(595),
(593),
(591),
(590),
(588),
(587),
(585),
(583),
(582),
(580),
(578),
(577),
(575),
(573),
(572),
(570),
(568),
(567),
(565),
(563),
(562),
(560),
(558),
(557),
(555),
(553),
(552),
(550),
(548),
(547),
(545),
(543),
(542),
(540),
(539),
(537),
(535),
(534),
(532),
(530),
(529),
(527),
(525),
(524),
(522),
(520),
(519),
(517),
(515),
(514),
(512),
(510),
(509),
(507),
(505),
(504),
(502),
(500),
(499),
(497),
(495),
(494),
(492),
(491),
(489),
(487),
(486),
(484),
(482),
(481),
(479),
(477),
(476),
(474),
(472),
(471),
(469),
(467),
(466),
(464),
(462),
(461),
(459),
(457),
(456),
(454),
(452),
(451),
(449),
(447),
(446),
(444),
(443),
(441),
(439),
(438),
(436),
(434),
(433),
(431),
(429),
(428),
(426),
(424),
(423),
(421),
(419),
(418),
(416),
(414),
(413),
(411),
(409),
(408),
(406),
(404),
(403),
(401),
(399),
(398),
(396),
(395),
(393),
(391),
(390),
(388),
(386),
(385),
(383),
(381),
(380),
(378),
(376),
(375),
(373),
(371),
(370),
(368),
(366),
(365),
(363),
(361),
(360),
(358),
(356),
(355),
(353),
(352),
(350),
(348),
(347),
(345),
(343),
(342),
(340),
(338),
(337),
(335),
(333),
(332),
(330),
(328),
(327),
(325),
(323),
(322),
(320),
(318),
(317),
(315),
(313),
(312),
(310),
(308),
(307),
(305),
(304),
(302),
(300),
(299),
(297),
(295),
(294),
(292),
(290),
(289),
(287),
(285),
(284),
(282),
(280),
(279),
(277),
(275),
(274),
(272),
(270),
(269),
(267),
(265),
(264),
(262),
(260),
(259),
(257),
(256),
(254),
(252),
(251),
(249),
(247),
(246),
(244),
(242),
(241),
(239),
(237),
(236),
(234),
(232),
(231),
(229),
(227),
(226),
(224),
(222),
(221),
(219),
(217),
(216),
(214),
(212),
(211),
(209),
(208),
(206),
(204),
(203),
(201),
(199),
(198),
(196),
(194),
(193),
(191),
(189),
(188),
(186),
(184),
(183),
(181),
(179),
(178),
(176),
(174),
(173),
(171),
(169),
(168),
(166),
(164),
(163),
(161),
(160),
(158),
(156),
(155),
(153),
(151),
(150),
(148),
(146),
(145),
(143),
(141),
(140),
(138),
(136),
(135),
(133),
(131),
(130),
(128),
(126),
(125),
(123),
(121),
(120),
(118),
(117),
(115),
(113),
(112),
(110),
(108),
(107),
(105),
(103),
(102),
(100),
(98),
(97),
(95),
(93),
(92),
(90),
(88),
(87),
(85),
(83),
(82),
(80),
(78),
(77),
(75),
(73),
(72),
(70),
(69),
(67),
(65),
(64),
(62),
(60),
(59),
(57),
(55),
(54),
(52),
(50),
(49),
(47),
(45),
(44),
(42),
(40),
(39),
(37),
(35),
(34),
(32),
(30),
(29),
(27),
(25),
(24),
(22),
(21),
(19),
(17),
(16),
(14),
(12),
(11),
(9),
(7),
(6),
(4),
(2),
(1),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095),
(4095)
);


begin
    -- This is the only statement required. It looks up the converted value of 
	-- the voltage input (in mV) in the v2d_LUT look-up table, and outputs the 
	-- distance (in 10^-4 m) in std_logic_vector format.
		yeet : process(index)
	begin
	if(rising_edge(clk)) then
		if(index < 0) then
			Amplitude <= 4095;
		elsif (index > 4095) then
			Amplitude <= 4095;
		else
			Amplitude <= BuzzAmps(index);
		end if;
	end if;
	end process;
--   distance <= std_logic_vector(to_unsigned(v2d_LUTshort(to_integer(unsigned(voltage))),distance'length));
--   distance <= std_logic_vector(to_unsigned(v2d_LUT(to_integer(unsigned(voltage))),distance'length));

end behavior;
