
-- In this example, we're going to map voltage to distance, using a linear 
-- approximation, according to the Sharp GP2Y0A41SK0F datasheet page 4, or 
-- Lab 3 handout page 5. 
-- 
-- The relevant points we will select are:
-- 2.750 V is  4.00 cm (or 2750 mV and  40.0 mm)
-- 0.400 V is 33.00 cm (or  400 mV and 330.0 mm)
-- 
-- Mapping to the scales in our system
-- 2750 (mV) should map to  400 (10^-4 m)
--  400 (mV) should map to 3300 (10^-4 m)
-- and developing a linear equation, we find:
--
-- Distance = -2900/2350 * Voltage + 3793.617
-- Note this code implements linear function, you must map to the 
-- NON-linear relationship in the datasheet. This code is only provided 
-- for reference to help get you started.

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY BuzzFreq_Lookup IS
   PORT(
      clk            :  IN    STD_LOGIC;                                
      reset          :  IN    STD_LOGIC;                                
      index      	 :  IN    integer;                           
      Increment     :  OUT   integer
		);
END BuzzFreq_Lookup;

ARCHITECTURE behavior OF BuzzFreq_Lookup IS

type array_1d is array (0 to 4095) of Integer;

constant Increments : array_1d := (						
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(56951266),
(56950479),
(56949692),
(56948904),
(56948117),
(56947329),
(56946542),
(56945754),
(56944967),
(56944180),
(56943392),
(56942605),
(56941817),
(56941030),
(56940243),
(56939455),
(56938668),
(56937880),
(56937093),
(56936306),
(56935518),
(56934731),
(56933943),
(56933156),
(56932368),
(56931581),
(56930794),
(56930006),
(56929219),
(56928431),
(56927644),
(56926857),
(56926069),
(56925282),
(56924494),
(56923707),
(56922920),
(56922132),
(56921345),
(56920557),
(56919770),
(56918983),
(56918195),
(56917408),
(56916620),
(56915833),
(56915045),
(56914258),
(56913471),
(56912683),
(56911896),
(56911108),
(56910321),
(56909534),
(56908746),
(56907959),
(56907171),
(56906384),
(56905597),
(56904809),
(56904022),
(56903234),
(56902447),
(56901659),
(56900872),
(56900085),
(56899297),
(56898510),
(56897722),
(56896935),
(56896148),
(56895360),
(56894573),
(56893785),
(56892998),
(56892211),
(56891423),
(56890636),
(56889848),
(56889061),
(56888273),
(56887486),
(56886699),
(56885911),
(56885124),
(56884336),
(56883549),
(56882762),
(56881974),
(56881187),
(56880399),
(56879612),
(56878825),
(56878037),
(56877250),
(56876462),
(56875675),
(56874888),
(56874100),
(56873313),
(56872525),
(56871738),
(56870950),
(56870163),
(56869376),
(56868588),
(56867801),
(56867013),
(56866226),
(56865439),
(56864651),
(56863864),
(56863076),
(56862289),
(56861502),
(56860714),
(56859927),
(56859139),
(56858352),
(56857564),
(56856777),
(56855990),
(56855202),
(56854415),
(56853627),
(56852840),
(56852053),
(56851265),
(56850478),
(56849690),
(56848903),
(56848116),
(56847328),
(56846541),
(56845753),
(56844966),
(56844178),
(56843391),
(56842604),
(56841816),
(56841029),
(56840241),
(56839454),
(56838667),
(56837879),
(56837092),
(56836304),
(56835517),
(56834730),
(56833942),
(56833155),
(56832367),
(56831580),
(56830793),
(56830005),
(56829218),
(56828430),
(56827643),
(56826855),
(56826068),
(56825281),
(56824493),
(56823706),
(56822918),
(56822131),
(56821344),
(56820556),
(56819769),
(56818981),
(56818194),
(56817407),
(56816619),
(56815832),
(56815044),
(56814257),
(56813469),
(56812682),
(56811895),
(56811107),
(56810320),
(56809532),
(56808745),
(56807958),
(56807170),
(56806383),
(56805595),
(56804808),
(56804021),
(56803233),
(56802446),
(56801658),
(56800871),
(56800083),
(56799296),
(56798509),
(56797721),
(56796934),
(56796146),
(56795359),
(56794572),
(56793784),
(56792997),
(56792209),
(56791422),
(56790635),
(56789847),
(56789060),
(56788272),
(56787485),
(56786698),
(56785910),
(56785123),
(56784335),
(56783548),
(56782760),
(56781973),
(56781186),
(56780398),
(56779611),
(56778823),
(56778036),
(56777249),
(56776461),
(56775674),
(56774886),
(56774099),
(56773312),
(56772524),
(56771737),
(56770949),
(56770162),
(56769374),
(56768587),
(56767800),
(56767012),
(56766225),
(56765437),
(56764650),
(56763863),
(56763075),
(56762288),
(56761500),
(56760713),
(56759926),
(56759138),
(56758351),
(56757563),
(56756776),
(56755988),
(56755201),
(56754414),
(56753626),
(56752839),
(56752051),
(56751264),
(56750477),
(56749689),
(56748902),
(56748114),
(56747327),
(56746540),
(56745752),
(56744965),
(56744177),
(56743390),
(56742603),
(56741815),
(56741028),
(56740240),
(56739453),
(56738665),
(56737878),
(56737091),
(56736303),
(56735516),
(56734728),
(56733941),
(56733154),
(56732366),
(56731579),
(56730791),
(56730004),
(56729217),
(56728429),
(56727642),
(56726854),
(56726067),
(56725279),
(56724492),
(56723705),
(56722917),
(56722130),
(56721342),
(56720555),
(56719768),
(56718980),
(56718193),
(56717405),
(56716618),
(56715831),
(56715043),
(56714256),
(56713468),
(56712681),
(56711894),
(56711106),
(56710319),
(56709531),
(56708744),
(56707956),
(56707169),
(56706382),
(56705594),
(56704807),
(56704019),
(56703232),
(56702445),
(56701657),
(56700870),
(56700082),
(56699295),
(56698508),
(56697720),
(56696933),
(56696145),
(56695358),
(56694570),
(56693783),
(56692996),
(56692208),
(56691421),
(56690633),
(56689846),
(56689059),
(56688271),
(56687484),
(56686696),
(56685909),
(56685122),
(56684334),
(56683547),
(56682759),
(56681972),
(56681184),
(56680397),
(56679610),
(56678822),
(56678035),
(56677247),
(56676460),
(56675673),
(56674885),
(56674098),
(56673310),
(56672523),
(56671736),
(56670948),
(56670161),
(56669373),
(56668586),
(56667799),
(56667011),
(56666224),
(56665436),
(56664649),
(56663861),
(56663074),
(56662287),
(56661499),
(56660712),
(56659924),
(56659137),
(56658350),
(56657562),
(56656775),
(56655987),
(56655200),
(56654413),
(56653625),
(56652838),
(56652050),
(56651263),
(56650475),
(56649688),
(56648901),
(56648113),
(56647326),
(56646538),
(56645751),
(56644964),
(56644176),
(56643389),
(56642601),
(56641814),
(56641027),
(56640239),
(56639452),
(56638664),
(56637877),
(56637089),
(56636302),
(56635515),
(56634727),
(56633940),
(56633152),
(56632365),
(56631578),
(56630790),
(56630003),
(56629215),
(56628428),
(56627641),
(56626853),
(56626066),
(56625278),
(56624491),
(56623704),
(56622916),
(56622129),
(56621341),
(56620554),
(56619766),
(56618979),
(56618192),
(56617404),
(56616617),
(56615829),
(56615042),
(56614255),
(56613467),
(56612680),
(56611892),
(56611105),
(56610318),
(56609530),
(56608743),
(56607955),
(56607168),
(56606380),
(56605593),
(56604806),
(56604018),
(56603231),
(56602443),
(56601656),
(56600869),
(56600081),
(56599294),
(56598506),
(56597719),
(56596932),
(56596144),
(56595357),
(56594569),
(56593782),
(56592994),
(56592207),
(56591420),
(56590632),
(56589845),
(56589057),
(56588270),
(56587483),
(56586695),
(56585908),
(56585120),
(56584333),
(56583546),
(56582758),
(56581971),
(56581183),
(56580396),
(56579609),
(56578821),
(56578034),
(56577246),
(56576459),
(56575671),
(56574884),
(56574097),
(56573309),
(56572522),
(56571734),
(56570947),
(56570160),
(56569372),
(56568585),
(56567797),
(56567010),
(56566223),
(56565435),
(56564648),
(56563860),
(56563073),
(56562285),
(56561498),
(56560711),
(56559923),
(56559136),
(56558348),
(56557561),
(56556774),
(56555986),
(56555199),
(56554411),
(56553624),
(56552837),
(56552049),
(56551262),
(56550474),
(56549687),
(56548899),
(56548112),
(56547325),
(56546537),
(56545750),
(56544962),
(56544175),
(56543388),
(56542600),
(56541813),
(56541025),
(56540238),
(56539451),
(56538663),
(56537876),
(56537088),
(56536301),
(56535514),
(56534726),
(56533939),
(56533151),
(56532364),
(56531576),
(56530789),
(56530002),
(56529214),
(56528427),
(56527639),
(56526852),
(56526065),
(56525277),
(56524490),
(56523702),
(56522915),
(56522128),
(56521340),
(56520553),
(56519765),
(56518978),
(56518190),
(56517403),
(56516616),
(56515828),
(56515041),
(56514253),
(56513466),
(56512679),
(56511891),
(56511104),
(56510316),
(56509529),
(56508742),
(56507954),
(56507167),
(56506379),
(56505592),
(56504804),
(56504017),
(56503230),
(56502442),
(56501655),
(56500867),
(56500080),
(56499293),
(56498505),
(56497718),
(56496930),
(56496143),
(56495356),
(56494568),
(56493781),
(56492993),
(56492206),
(56491419),
(56490631),
(56489844),
(56489056),
(56488269),
(56487481),
(56486694),
(56485907),
(56485119),
(56484332),
(56483544),
(56482757),
(56481970),
(56481182),
(56480395),
(56479607),
(56478820),
(56478033),
(56477245),
(56476458),
(56475670),
(56474883),
(56474095),
(56473308),
(56472521),
(56471733),
(56470946),
(56470158),
(56469371),
(56468584),
(56467796),
(56467009),
(56466221),
(56465434),
(56464647),
(56463859),
(56463072),
(56462284),
(56461497),
(56460709),
(56459922),
(56459135),
(56458347),
(56457560),
(56456772),
(56455985),
(56455198),
(56454410),
(56453623),
(56452835),
(56452048),
(56451261),
(56450473),
(56449686),
(56448898),
(56448111),
(56447324),
(56446536),
(56445749),
(56444961),
(56444174),
(56443386),
(56442599),
(56441812),
(56441024),
(56440237),
(56439449),
(56438662),
(56437875),
(56437087),
(56436300),
(56435512),
(56434725),
(56433938),
(56433150),
(56432363),
(56431575),
(56430788),
(56430000),
(56429213),
(56428426),
(56427638),
(56426851),
(56426063),
(56425276),
(56424489),
(56423701),
(56422914),
(56422126),
(56421339),
(56420552),
(56419764),
(56418977),
(56418189),
(56417402),
(56416614),
(56415827),
(56415040),
(56414252),
(56413465),
(56412677),
(56411890),
(56411103),
(56410315),
(56409528),
(56408740),
(56407953),
(56407166),
(56406378),
(56405591),
(56404803),
(56404016),
(56403229),
(56402441),
(56401654),
(56400866),
(56400079),
(56399291),
(56398504),
(56397717),
(56396929),
(56396142),
(56395354),
(56394567),
(56393780),
(56392992),
(56392205),
(56391417),
(56390630),
(56389843),
(56389055),
(56388268),
(56387480),
(56386693),
(56385905),
(56385118),
(56384331),
(56383543),
(56382756),
(56381968),
(56381181),
(56380394),
(56379606),
(56378819),
(56378031),
(56377244),
(56376457),
(56375669),
(56374882),
(56374094),
(56373307),
(56372520),
(56371732),
(56370945),
(56370157),
(56369370),
(56368582),
(56367795),
(56367008),
(56366220),
(56365433),
(56364645),
(56363858),
(56363071),
(56362283),
(56361496),
(56360708),
(56359921),
(56359134),
(56358346),
(56357559),
(56356771),
(56355984),
(56355196),
(56354409),
(56353622),
(56352834),
(56352047),
(56351259),
(56350472),
(56349685),
(56348897),
(56348110),
(56347322),
(56346535),
(56345748),
(56344960),
(56344173),
(56343385),
(56342598),
(56341810),
(56341023),
(56340236),
(56339448),
(56338661),
(56337873),
(56337086),
(56336299),
(56335511),
(56334724),
(56333936),
(56333149),
(56332362),
(56331574),
(56330787),
(56329999),
(56329212),
(56328425),
(56327637),
(56326850),
(56326062),
(56325275),
(56324487),
(56323700),
(56322913),
(56322125),
(56321338),
(56320550),
(56319763),
(56318976),
(56318188),
(56317401),
(56316613),
(56315826),
(56315039),
(56314251),
(56313464),
(56312676),
(56311889),
(56311101),
(56310314),
(56309527),
(56308739),
(56307952),
(56307164),
(56306377),
(56305590),
(56304802),
(56304015),
(56303227),
(56302440),
(56301653),
(56300865),
(56300078),
(56299290),
(56298503),
(56297715),
(56296928),
(56296141),
(56295353),
(56294566),
(56293778),
(56292991),
(56292204),
(56291416),
(56290629),
(56289841),
(56289054),
(56288267),
(56287479),
(56286692),
(56285904),
(56285117),
(56284330),
(56283542),
(56282755),
(56281967),
(56281180),
(56280392),
(56279605),
(56278818),
(56278030),
(56277243),
(56276455),
(56275668),
(56274881),
(56274093),
(56273306),
(56272518),
(56271731),
(56270944),
(56270156),
(56269369),
(56268581),
(56267794),
(56267006),
(56266219),
(56265432),
(56264644),
(56263857),
(56263069),
(56262282),
(56261495),
(56260707),
(56259920),
(56259132),
(56258345),
(56257558),
(56256770),
(56255983),
(56255195),
(56254408),
(56253620),
(56252833),
(56252046),
(56251258),
(56250471),
(56249683),
(56248896),
(56248109),
(56247321),
(56246534),
(56245746),
(56244959),
(56244172),
(56243384),
(56242597),
(56241809),
(56241022),
(56240235),
(56239447),
(56238660),
(56237872),
(56237085),
(56236297),
(56235510),
(56234723),
(56233935),
(56233148),
(56232360),
(56231573),
(56230786),
(56229998),
(56229211),
(56228423),
(56227636),
(56226849),
(56226061),
(56225274),
(56224486),
(56223699),
(56222911),
(56222124),
(56221337),
(56220549),
(56219762),
(56218974),
(56218187),
(56217400),
(56216612),
(56215825),
(56215037),
(56214250),
(56213463),
(56212675),
(56211888),
(56211100),
(56210313),
(56209525),
(56208738),
(56207951),
(56207163),
(56206376),
(56205588),
(56204801),
(56204014),
(56203226),
(56202439),
(56201651),
(56200864),
(56200077),
(56199289),
(56198502),
(56197714),
(56196927),
(56196140),
(56195352),
(56194565),
(56193777),
(56192990),
(56192202),
(56191415),
(56190628),
(56189840),
(56189053),
(56188265),
(56187478),
(56186691),
(56185903),
(56185116),
(56184328),
(56183541),
(56182754),
(56181966),
(56181179),
(56180391),
(56179604),
(56178816),
(56178029),
(56177242),
(56176454),
(56175667),
(56174879),
(56174092),
(56173305),
(56172517),
(56171730),
(56170942),
(56170155),
(56169368),
(56168580),
(56167793),
(56167005),
(56166218),
(56165430),
(56164643),
(56163856),
(56163068),
(56162281),
(56161493),
(56160706),
(56159919),
(56159131),
(56158344),
(56157556),
(56156769),
(56155982),
(56155194),
(56154407),
(56153619),
(56152832),
(56152045),
(56151257),
(56150470),
(56149682),
(56148895),
(56148107),
(56147320),
(56146533),
(56145745),
(56144958),
(56144170),
(56143383),
(56142596),
(56141808),
(56141021),
(56140233),
(56139446),
(56138659),
(56137871),
(56137084),
(56136296),
(56135509),
(56134721),
(56133934),
(56133147),
(56132359),
(56131572),
(56130784),
(56129997),
(56129210),
(56128422),
(56127635),
(56126847),
(56126060),
(56125273),
(56124485),
(56123698),
(56122910),
(56122123),
(56121335),
(56120548),
(56119761),
(56118973),
(56118186),
(56117398),
(56116611),
(56115824),
(56115036),
(56114249),
(56113461),
(56112674),
(56111887),
(56111099),
(56110312),
(56109524),
(56108737),
(56107950),
(56107162),
(56106375),
(56105587),
(56104800),
(56104012),
(56103225),
(56102438),
(56101650),
(56100863),
(56100075),
(56099288),
(56098501),
(56097713),
(56096926),
(56096138),
(56095351),
(56094564),
(56093776),
(56092989),
(56092201),
(56091414),
(56090626),
(56089839),
(56089052),
(56088264),
(56087477),
(56086689),
(56085902),
(56085115),
(56084327),
(56083540),
(56082752),
(56081965),
(56081178),
(56080390),
(56079603),
(56078815),
(56078028),
(56077241),
(56076453),
(56075666),
(56074878),
(56074091),
(56073303),
(56072516),
(56071729),
(56070941),
(56070154),
(56069366),
(56068579),
(56067792),
(56067004),
(56066217),
(56065429),
(56064642),
(56063855),
(56063067),
(56062280),
(56061492),
(56060705),
(56059917),
(56059130),
(56058343),
(56057555),
(56056768),
(56055980),
(56055193),
(56054406),
(56053618),
(56052831),
(56052043),
(56051256),
(56050469),
(56049681),
(56048894),
(56048106),
(56047319),
(56046531),
(56045744),
(56044957),
(56044169),
(56043382),
(56042594),
(56041807),
(56041020),
(56040232),
(56039445),
(56038657),
(56037870),
(56037083),
(56036295),
(56035508),
(56034720),
(56033933),
(56033146),
(56032358),
(56031571),
(56030783),
(56029996),
(56029208),
(56028421),
(56027634),
(56026846),
(56026059),
(56025271),
(56024484),
(56023697),
(56022909),
(56022122),
(56021334),
(56020547),
(56019760),
(56018972),
(56018185),
(56017397),
(56016610),
(56015822),
(56015035),
(56014248),
(56013460),
(56012673),
(56011885),
(56011098),
(56010311),
(56009523),
(56008736),
(56007948),
(56007161),
(56006374),
(56005586),
(56004799),
(56004011),
(56003224),
(56002436),
(56001649),
(56000862),
(56000074),
(55999287),
(55998499),
(55997712),
(55996925),
(55996137),
(55995350),
(55994562),
(55993775),
(55992988),
(55992200),
(55991413),
(55990625),
(55989838),
(55989051),
(55988263),
(55987476),
(55986688),
(55985901),
(55985113),
(55984326),
(55983539),
(55982751),
(55981964),
(55981176),
(55980389),
(55979602),
(55978814),
(55978027),
(55977239),
(55976452),
(55975665),
(55974877),
(55974090),
(55973302),
(55972515),
(55971727),
(55970940),
(55970153),
(55969365),
(55968578),
(55967790),
(55967003),
(55966216),
(55965428),
(55964641),
(55963853),
(55963066),
(55962279),
(55961491),
(55960704),
(55959916),
(55959129),
(55958341),
(55957554),
(55956767),
(55955979),
(55955192),
(55954404),
(55953617),
(55952830),
(55952042),
(55951255),
(55950467),
(55949680),
(55948893),
(55948105),
(55947318),
(55946530),
(55945743),
(55944956),
(55944168),
(55943381),
(55942593),
(55941806),
(55941018),
(55940231),
(55939444),
(55938656),
(55937869),
(55937081),
(55936294),
(55935507),
(55934719),
(55933932),
(55933144),
(55932357),
(55931570),
(55930782),
(55929995),
(55929207),
(55928420),
(55927632),
(55926845),
(55926058),
(55925270),
(55924483),
(55923695),
(55922908),
(55922121),
(55921333),
(55920546),
(55919758),
(55918971),
(55918184),
(55917396),
(55916609),
(55915821),
(55915034),
(55914246),
(55913459),
(55912672),
(55911884),
(55911097),
(55910309),
(55909522),
(55908735),
(55907947),
(55907160),
(55906372),
(55905585),
(55904798),
(55904010),
(55903223),
(55902435),
(55901648),
(55900861),
(55900073),
(55899286),
(55898498),
(55897711),
(55896923),
(55896136),
(55895349),
(55894561),
(55893774),
(55892986),
(55892199),
(55891412),
(55890624),
(55889837),
(55889049),
(55888262),
(55887475),
(55886687),
(55885900),
(55885112),
(55884325),
(55883537),
(55882750),
(55881963),
(55881175),
(55880388),
(55879600),
(55878813),
(55878026),
(55877238),
(55876451),
(55875663),
(55874876),
(55874089),
(55873301),
(55872514),
(55871726),
(55870939),
(55870151),
(55869364),
(55868577),
(55867789),
(55867002),
(55866214),
(55865427),
(55864640),
(55863852),
(55863065),
(55862277),
(55861490),
(55860703),
(55859915),
(55859128),
(55858340),
(55857553),
(55856766),
(55855978),
(55855191),
(55854403),
(55853616),
(55852828),
(55852041),
(55851254),
(55850466),
(55849679),
(55848891),
(55848104),
(55847317),
(55846529),
(55845742),
(55844954),
(55844167),
(55843380),
(55842592),
(55841805),
(55841017),
(55840230),
(55839442),
(55838655),
(55837868),
(55837080),
(55836293),
(55835505),
(55834718),
(55833931),
(55833143),
(55832356),
(55831568),
(55830781),
(55829994),
(55829206),
(55828419),
(55827631),
(55826844),
(55826056),
(55825269),
(55824482),
(55823694),
(55822907),
(55822119),
(55821332),
(55820545),
(55819757),
(55818970),
(55818182),
(55817395),
(55816608),
(55815820),
(55815033),
(55814245),
(55813458),
(55812671),
(55811883),
(55811096),
(55810308),
(55809521),
(55808733),
(55807946),
(55807159),
(55806371),
(55805584),
(55804796),
(55804009),
(55803222),
(55802434),
(55801647),
(55800859),
(55800072),
(55799285),
(55798497),
(55797710),
(55796922),
(55796135),
(55795347),
(55794560),
(55793773),
(55792985),
(55792198),
(55791410),
(55790623),
(55789836),
(55789048),
(55788261),
(55787473),
(55786686),
(55785899),
(55785111),
(55784324),
(55783536),
(55782749),
(55781961),
(55781174),
(55780387),
(55779599),
(55778812),
(55778024),
(55777237),
(55776450),
(55775662),
(55774875),
(55774087),
(55773300),
(55772513),
(55771725),
(55770938),
(55770150),
(55769363),
(55768576),
(55767788),
(55767001),
(55766213),
(55765426),
(55764638),
(55763851),
(55763064),
(55762276),
(55761489),
(55760701),
(55759914),
(55759127),
(55758339),
(55757552),
(55756764),
(55755977),
(55755190),
(55754402),
(55753615),
(55752827),
(55752040),
(55751252),
(55750465),
(55749678),
(55748890),
(55748103),
(55747315),
(55746528),
(55745741),
(55744953),
(55744166),
(55743378),
(55742591),
(55741804),
(55741016),
(55740229),
(55739441),
(55738654),
(55737867),
(55737079),
(55736292),
(55735504),
(55734717),
(55733929),
(55733142),
(55732355),
(55731567),
(55730780),
(55729992),
(55729205),
(55728418),
(55727630),
(55726843),
(55726055),
(55725268),
(55724481),
(55723693),
(55722906),
(55722118),
(55721331),
(55720543),
(55719756),
(55718969),
(55718181),
(55717394),
(55716606),
(55715819),
(55715032),
(55714244),
(55713457),
(55712669),
(55711882),
(55711095),
(55710307),
(55709520),
(55708732),
(55707945),
(55707157),
(55706370),
(55705583),
(55704795),
(55704008),
(55703220),
(55702433),
(55701646),
(55700858),
(55700071),
(55699283),
(55698496),
(55697709),
(55696921),
(55696134),
(55695346),
(55694559),
(55693772),
(55692984),
(55692197),
(55691409),
(55690622),
(55689834),
(55689047),
(55688260),
(55687472),
(55686685),
(55685897),
(55685110),
(55684323),
(55683535),
(55682748),
(55681960),
(55681173),
(55680386),
(55679598),
(55678811),
(55678023),
(55677236),
(55676448),
(55675661),
(55674874),
(55674086),
(55673299),
(55672511),
(55671724),
(55670937),
(55670149),
(55669362),
(55668574),
(55667787),
(55667000),
(55666212),
(55665425),
(55664637),
(55663850),
(55663062),
(55662275),
(55661488),
(55660700),
(55659913),
(55659125),
(55658338),
(55657551),
(55656763),
(55655976),
(55655188),
(55654401),
(55653614),
(55652826),
(55652039),
(55651251),
(55650464),
(55649677),
(55648889),
(55648102),
(55647314),
(55646527),
(55645739),
(55644952),
(55644165),
(55643377),
(55642590),
(55641802),
(55641015),
(55640228),
(55639440),
(55638653),
(55637865),
(55637078),
(55636291),
(55635503),
(55634716),
(55633928),
(55633141),
(55632353),
(55631566),
(55630779),
(55629991),
(55629204),
(55628416),
(55627629),
(55626842),
(55626054),
(55625267),
(55624479),
(55623692),
(55622905),
(55622117),
(55621330),
(55620542),
(55619755),
(55618967),
(55618180),
(55617393),
(55616605),
(55615818),
(55615030),
(55614243),
(55613456),
(55612668),
(55611881),
(55611093),
(55610306),
(55609519),
(55608731),
(55607944),
(55607156),
(55606369),
(55605582),
(55604794),
(55604007),
(55603219),
(55602432),
(55601644),
(55600857),
(55600070),
(55599282),
(55598495),
(55597707),
(55596920),
(55596133),
(55595345),
(55594558),
(55593770),
(55592983),
(55592196),
(55591408),
(55590621),
(55589833),
(55589046),
(55588258),
(55587471),
(55586684),
(55585896),
(55585109),
(55584321),
(55583534),
(55582747),
(55581959),
(55581172),
(55580384),
(55579597),
(55578810),
(55578022),
(55577235),
(55576447),
(55575660),
(55574872),
(55574085),
(55573298),
(55572510),
(55571723),
(55570935),
(55570148),
(55569361),
(55568573),
(55567786),
(55566998),
(55566211),
(55565424),
(55564636),
(55563849),
(55563061),
(55562274),
(55561487),
(55560699),
(55559912),
(55559124),
(55558337),
(55557549),
(55556762),
(55555975),
(55555187),
(55554400),
(55553612),
(55552825),
(55552038),
(55551250),
(55550463),
(55549675),
(55548888),
(55548101),
(55547313),
(55546526),
(55545738),
(55544951),
(55544163),
(55543376),
(55542589),
(55541801),
(55541014),
(55540226),
(55539439),
(55538652),
(55537864),
(55537077),
(55536289),
(55535502),
(55534715),
(55533927),
(55533140),
(55532352),
(55531565),
(55530777),
(55529990),
(55529203),
(55528415),
(55527628),
(55526840),
(55526053),
(55525266),
(55524478),
(55523691),
(55522903),
(55522116),
(55521329),
(55520541),
(55519754),
(55518966),
(55518179),
(55517392),
(55516604),
(55515817),
(55515029),
(55514242),
(55513454),
(55512667),
(55511880),
(55511092),
(55510305),
(55509517),
(55508730),
(55507943),
(55507155),
(55506368),
(55505580),
(55504793),
(55504006),
(55503218),
(55502431),
(55501643),
(55500856),
(55500068),
(55499281),
(55498494),
(55497706),
(55496919),
(55496131),
(55495344),
(55494557),
(55493769),
(55492982),
(55492194),
(55491407),
(55490620),
(55489832),
(55489045),
(55488257),
(55487470),
(55486682),
(55485895),
(55485108),
(55484320),
(55483533),
(55482745),
(55481958),
(55481171),
(55480383),
(55479596),
(55478808),
(55478021),
(55477234),
(55476446),
(55475659),
(55474871),
(55474084),
(55473297),
(55472509),
(55471722),
(55470934),
(55470147),
(55469359),
(55468572),
(55467785),
(55466997),
(55466210),
(55465422),
(55464635),
(55463848),
(55463060),
(55462273),
(55461485),
(55460698),
(55459911),
(55459123),
(55458336),
(55457548),
(55456761),
(55455973),
(55455186),
(55454399),
(55453611),
(55452824),
(55452036),
(55451249),
(55450462),
(55449674),
(55448887),
(55448099),
(55447312),
(55446525),
(55445737),
(55444950),
(55444162),
(55443375),
(55442587),
(55441800),
(55441013),
(55440225),
(55439438),
(55438650),
(55437863),
(55437076),
(55436288),
(55435501),
(55434713),
(55433926),
(55433139),
(55432351),
(55431564),
(55430776),
(55429989),
(55429202),
(55428414),
(55427627),
(55426839),
(55426052),
(55425264),
(55424477),
(55423690),
(55422902),
(55422115),
(55421327),
(55420540),
(55419753),
(55418965),
(55418178),
(55417390),
(55416603),
(55415816),
(55415028),
(55414241),
(55413453),
(55412666),
(55411878),
(55411091),
(55410304),
(55409516),
(55408729),
(55407941),
(55407154),
(55406367),
(55405579),
(55404792),
(55404004),
(55403217),
(55402430),
(55401642),
(55400855),
(55400067),
(55399280),
(55398493),
(55397705),
(55396918),
(55396130),
(55395343),
(55394555),
(55393768),
(55392981),
(55392193),
(55391406),
(55390618),
(55389831),
(55389044),
(55388256),
(55387469),
(55386681),
(55385894),
(55385107),
(55384319),
(55383532),
(55382744),
(55381957),
(55381169),
(55380382),
(55379595),
(55378807),
(55378020),
(55377232),
(55376445),
(55375658),
(55374870),
(55374083),
(55373295),
(55372508),
(55371721),
(55370933),
(55370146),
(55369358),
(55368571),
(55367783),
(55366996),
(55366209),
(55365421),
(55364634),
(55363846),
(55363059),
(55362272),
(55361484),
(55360697),
(55359909),
(55359122),
(55358335),
(55357547),
(55356760),
(55355972),
(55355185),
(55354398),
(55353610),
(55352823),
(55352035),
(55351248),
(55350460),
(55349673),
(55348886),
(55348098),
(55347311),
(55346523),
(55345736),
(55344949),
(55344161),
(55343374),
(55342586),
(55341799),
(55341012),
(55340224),
(55339437),
(55338649),
(55337862),
(55337074),
(55336287),
(55335500),
(55334712),
(55333925),
(55333137),
(55332350),
(55331563),
(55330775),
(55329988),
(55329200),
(55328413),
(55327626),
(55326838),
(55326051),
(55325263),
(55324476),
(55323688),
(55322901),
(55322114),
(55321326),
(55320539),
(55319751),
(55318964),
(55318177),
(55317389),
(55316602),
(55315814),
(55315027),
(55314240),
(55313452),
(55312665),
(55311877),
(55311090),
(55310303),
(55309515),
(55308728),
(55307940),
(55307153),
(55306365),
(55305578),
(55304791),
(55304003),
(55303216),
(55302428),
(55301641),
(55300854),
(55300066),
(55299279),
(55298491),
(55297704),
(55296917),
(55296129),
(55295342),
(55294554),
(55293767),
(55292979),
(55292192),
(55291405),
(55290617),
(55289830),
(55289042),
(55288255),
(55287468),
(55286680),
(55285893),
(55285105),
(55284318),
(55283531),
(55282743),
(55281956),
(55281168),
(55280381),
(55279593),
(55278806),
(55278019),
(55277231),
(55276444),
(55275656),
(55274869),
(55274082),
(55273294),
(55272507),
(55271719),
(55270932),
(55270145),
(55269357),
(55268570),
(55267782),
(55266995),
(55266208),
(55265420),
(55264633),
(55263845),
(55263058),
(55262270),
(55261483),
(55260696),
(55259908),
(55259121),
(55258333),
(55257546),
(55256759),
(55255971),
(55255184),
(55254396),
(55253609),
(55252822),
(55252034),
(55251247),
(55250459),
(55249672),
(55248884),
(55248097),
(55247310),
(55246522),
(55245735),
(55244947),
(55244160),
(55243373),
(55242585),
(55241798),
(55241010),
(55240223),
(55239436),
(55238648),
(55237861),
(55237073),
(55236286),
(55235498),
(55234711),
(55233924),
(55233136),
(55232349),
(55231561),
(55230774),
(55229987),
(55229199),
(55228412),
(55227624),
(55226837),
(55226050),
(55225262),
(55224475),
(55223687),
(55222900),
(55222113),
(55221325),
(55220538),
(55219750),
(55218963),
(55218175),
(55217388),
(55216601),
(55215813),
(55215026),
(55214238),
(55213451),
(55212664),
(55211876),
(55211089),
(55210301),
(55209514),
(55208727),
(55207939),
(55207152),
(55206364),
(55205577),
(55204789),
(55204002),
(55203215),
(55202427),
(55201640),
(55200852),
(55200065),
(55199278),
(55198490),
(55197703),
(55196915),
(55196128),
(55195341),
(55194553),
(55193766),
(55192978),
(55192191),
(55191403),
(55190616),
(55189829),
(55189041),
(55188254),
(55187466),
(55186679),
(55185892),
(55185104),
(55184317),
(55183529),
(55182742),
(55181955),
(55181167),
(55180380),
(55179592),
(55178805),
(55178018),
(55177230),
(55176443),
(55175655),
(55174868),
(55174080),
(55173293),
(55172506),
(55171718),
(55170931),
(55170143),
(55169356),
(55168569),
(55167781),
(55166994),
(55166206),
(55165419),
(55164632),
(55163844),
(55163057),
(55162269),
(55161482),
(55160694),
(55159907),
(55159120),
(55158332),
(55157545),
(55156757),
(55155970),
(55155183),
(55154395),
(55153608),
(55152820),
(55152033),
(55151246),
(55150458),
(55149671),
(55148883),
(55148096),
(55147308),
(55146521),
(55145734),
(55144946),
(55144159),
(55143371),
(55142584),
(55141797),
(55141009),
(55140222),
(55139434),
(55138647),
(55137860),
(55137072),
(55136285),
(55135497),
(55134710),
(55133923),
(55133135),
(55132348),
(55131560),
(55130773),
(55129985),
(55129198),
(55128411),
(55127623),
(55126836),
(55126048),
(55125261),
(55124474),
(55123686),
(55122899),
(55122111),
(55121324),
(55120537),
(55119749),
(55118962),
(55118174),
(55117387),
(55116599),
(55115812),
(55115025),
(55114237),
(55113450),
(55112662),
(55111875),
(55111088),
(55110300),
(55109513),
(55108725),
(55107938),
(55107151),
(55106363),
(55105576),
(55104788),
(55104001),
(55103214),
(55102426),
(55101639),
(55100851),
(55100064),
(55099276),
(55098489),
(55097702),
(55096914),
(55096127),
(55095339),
(55094552),
(55093765),
(55092977),
(55092190),
(55091402),
(55090615),
(55089828),
(55089040),
(55088253),
(55087465),
(55086678),
(55085890),
(55085103),
(55084316),
(55083528),
(55082741),
(55081953),
(55081166),
(55080379),
(55079591),
(55078804),
(55078016),
(55077229),
(55076442),
(55075654),
(55074867),
(55074079),
(55073292),
(55072504),
(55071717),
(55070930),
(55070142),
(55069355),
(55068567),
(55067780),
(55066993),
(55066205),
(55065418),
(55064630),
(55063843),
(55063056),
(55062268),
(55061481),
(55060693),
(55059906),
(55059119),
(55058331),
(55057544),
(55056756),
(55055969),
(55055181),
(55054394),
(55053607),
(55052819),
(55052032),
(55051244),
(55050457),
(55049670),
(55048882),
(55048095),
(55047307),
(55046520),
(55045733),
(55044945),
(55044158),
(55043370),
(55042583),
(55041795),
(55041008),
(55040221),
(55039433),
(55038646),
(55037858),
(55037071),
(55036284),
(55035496),
(55034709),
(55033921),
(55033134),
(55032347),
(55031559),
(55030772),
(55029984),
(55029197),
(55028409),
(55027622),
(55026835),
(55026047),
(55025260),
(55024472),
(55023685),
(55022898),
(55022110),
(55021323),
(55020535),
(55019748),
(55018961),
(55018173),
(55017386),
(55016598),
(55015811),
(55015024),
(55014236),
(55013449),
(55012661),
(55011874),
(55011086),
(55010299),
(55009512),
(55008724),
(55007937),
(55007149),
(55006362),
(55005575),
(55004787),
(55004000),
(55003212),
(55002425),
(55001638),
(55000850),
(55000063),
(54999275),
(54998488),
(54997700),
(54996913),
(54996126),
(54995338),
(54994551),
(54993763),
(54992976),
(54992189),
(54991401),
(54990614),
(54989826),
(54989039),
(54988252),
(54987464),
(54986677),
(54985889),
(54985102),
(54984314),
(54983527),
(54982740),
(54981952),
(54981165),
(54980377),
(54979590),
(54978803),
(54978015),
(54977228),
(54976440),
(54975653),
(54974866),
(54974078),
(54973291),
(54972503),
(54971716),
(54970929),
(54970141),
(54969354),
(54968566),
(54967779),
(54966991),
(54966204),
(54965417),
(54964629),
(54963842),
(54963054),
(54962267),
(54961480),
(54960692),
(54959905),
(54959117),
(54958330),
(54957543),
(54956755),
(54955968),
(54955180),
(54954393),
(54953605),
(54952818),
(54952031),
(54951243),
(54950456),
(54949668),
(54948881),
(54948094),
(54947306),
(54946519),
(54945731),
(54944944),
(54944157),
(54943369),
(54942582),
(54941794),
(54941007),
(54940219),
(54939432),
(54938645),
(54937857),
(54937070),
(54936282),
(54935495),
(54934708),
(54933920),
(54933133),
(54932345),
(54931558),
(54930771),
(54929983),
(54929196),
(54928408),
(54927621),
(54926834),
(54926046),
(54925259),
(54924471),
(54923684),
(54922896),
(54922109),
(54921322),
(54920534),
(54919747),
(54918959),
(54918172),
(54917385),
(54916597),
(54915810),
(54915022),
(54914235),
(54913448),
(54912660),
(54911873),
(54911085),
(54910298),
(54909510),
(54908723),
(54907936),
(54907148),
(54906361),
(54905573),
(54904786),
(54903999),
(54903211),
(54902424),
(54901636),
(54900849),
(54900062),
(54899274),
(54898487),
(54897699),
(54896912),
(54896124),
(54895337),
(54894550),
(54893762),
(54892975),
(54892187),
(54891400),
(54890613),
(54889825),
(54889038),
(54888250),
(54887463),
(54886676),
(54885888),
(54885101),
(54884313),
(54883526),
(54882739),
(54881951),
(54881164),
(54880376),
(54879589),
(54878801),
(54878014),
(54877227),
(54876439),
(54875652),
(54874864),
(54874077),
(54873290),
(54872502),
(54871715),
(54870927),
(54870140),
(54869353),
(54868565),
(54867778),
(54866990),
(54866203),
(54865415),
(54864628),
(54863841),
(54863053),
(54862266),
(54861478),
(54860691),
(54859904),
(54859116),
(54858329),
(54857541),
(54856754),
(54855967),
(54855179),
(54854392),
(54853604),
(54852817),
(54852029),
(54851242),
(54850455),
(54849667),
(54848880),
(54848092),
(54847305),
(54846518),
(54845730),
(54844943),
(54844155),
(54843368),
(54842581),
(54841793),
(54841006),
(54840218),
(54839431),
(54838644),
(54837856),
(54837069),
(54836281),
(54835494),
(54834706),
(54833919),
(54833132),
(54832344),
(54831557),
(54830769),
(54829982),
(54829195),
(54828407),
(54827620),
(54826832),
(54826045),
(54825258),
(54824470),
(54823683),
(54822895),
(54822108),
(54821320),
(54820533),
(54819746),
(54818958),
(54818171),
(54817383),
(54816596),
(54815809),
(54815021),
(54814234),
(54813446),
(54812659),
(54811872),
(54811084),
(54810297),
(54809509),
(54808722),
(54807934),
(54807147),
(54806360),
(54805572),
(54804785),
(54803997),
(54803210),
(54802423),
(54801635),
(54800848),
(54800060),
(54799273),
(54798486),
(54797698),
(54796911),
(54796123),
(54795336),
(54794549),
(54793761),
(54792974),
(54792186),
(54791399),
(54790611),
(54789824),
(54789037),
(54788249),
(54787462),
(54786674),
(54785887),
(54785100),
(54784312),
(54783525),
(54782737),
(54781950),
(54781163),
(54780375),
(54779588),
(54778800),
(54778013),
(54777225),
(54776438),
(54775651),
(54774863),
(54774076),
(54773288),
(54772501),
(54771714),
(54770926),
(54770139),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575),
(55834575)
);


begin
    -- This is the only statement required. It looks up the converted value of 
	-- the voltage input (in mV) in the v2d_LUT look-up table, and outputs the 
	-- distance (in 10^-4 m) in std_logic_vector format.
	yeet : process(index)
	begin
		if(index < 0) then
			Increment <= 55834575;
		elsif (index > 4095) then
			Increment <= 55834575;
		else
			Increment <= Increments(index);
		end if;
	end process;
--   distance <= std_logic_vector(to_unsigned(v2d_LUTshort(to_integer(unsigned(voltage))),distance'length));
--   distance <= std_logic_vector(to_unsigned(v2d_LUT(to_integer(unsigned(voltage))),distance'length));

end behavior;
